-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_727_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1061_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1011_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1061_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_1 : boolean;
  signal type_cast_538_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_1 : boolean;
  signal array_obj_ref_1362_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_req_0 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1029_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 : boolean;
  signal type_cast_1401_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_0 : boolean;
  signal addr_of_689_final_reg_ack_1 : boolean;
  signal type_cast_592_inst_ack_0 : boolean;
  signal type_cast_592_inst_req_0 : boolean;
  signal type_cast_538_inst_req_1 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_ack_1 : boolean;
  signal type_cast_709_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal if_stmt_632_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal WPIPE_Block0_start_973_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_0 : boolean;
  signal WPIPE_Block0_start_973_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_0 : boolean;
  signal ptr_deref_618_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 : boolean;
  signal type_cast_696_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_997_inst_ack_1 : boolean;
  signal type_cast_51_inst_req_0 : boolean;
  signal type_cast_51_inst_ack_0 : boolean;
  signal type_cast_51_inst_req_1 : boolean;
  signal type_cast_51_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1011_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1058_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1064_inst_req_1 : boolean;
  signal addr_of_689_final_reg_req_1 : boolean;
  signal WPIPE_Block1_start_1014_inst_req_1 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1011_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1014_inst_ack_1 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal type_cast_727_inst_req_1 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal type_cast_574_inst_ack_1 : boolean;
  signal type_cast_1371_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 : boolean;
  signal type_cast_574_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_997_inst_req_0 : boolean;
  signal if_stmt_632_branch_req_0 : boolean;
  signal WPIPE_Block0_start_982_inst_req_0 : boolean;
  signal array_obj_ref_688_index_offset_ack_1 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_req_1 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_982_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1079_inst_ack_0 : boolean;
  signal addr_of_689_final_reg_ack_0 : boolean;
  signal array_obj_ref_688_index_offset_req_1 : boolean;
  signal type_cast_101_inst_req_0 : boolean;
  signal type_cast_101_inst_ack_0 : boolean;
  signal type_cast_101_inst_req_1 : boolean;
  signal type_cast_101_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_973_inst_req_0 : boolean;
  signal type_cast_659_inst_ack_1 : boolean;
  signal type_cast_659_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 : boolean;
  signal type_cast_574_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 : boolean;
  signal type_cast_696_inst_ack_1 : boolean;
  signal type_cast_610_inst_ack_1 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1011_inst_req_1 : boolean;
  signal type_cast_574_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1051_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 : boolean;
  signal type_cast_696_inst_req_1 : boolean;
  signal addr_of_689_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 : boolean;
  signal type_cast_610_inst_req_1 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal array_obj_ref_688_index_offset_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal type_cast_659_inst_ack_0 : boolean;
  signal type_cast_1431_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_0 : boolean;
  signal type_cast_339_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_1 : boolean;
  signal type_cast_339_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_982_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_991_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_991_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_ack_1 : boolean;
  signal type_cast_138_inst_req_0 : boolean;
  signal ptr_deref_618_store_0_req_0 : boolean;
  signal type_cast_138_inst_ack_0 : boolean;
  signal array_obj_ref_688_index_offset_req_0 : boolean;
  signal type_cast_138_inst_req_1 : boolean;
  signal type_cast_138_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1079_inst_req_0 : boolean;
  signal type_cast_659_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1029_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 : boolean;
  signal type_cast_696_inst_req_0 : boolean;
  signal WPIPE_Block0_start_973_inst_req_1 : boolean;
  signal type_cast_151_inst_req_0 : boolean;
  signal type_cast_151_inst_ack_0 : boolean;
  signal type_cast_151_inst_req_1 : boolean;
  signal type_cast_151_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 : boolean;
  signal type_cast_163_inst_req_0 : boolean;
  signal type_cast_163_inst_ack_0 : boolean;
  signal type_cast_163_inst_req_1 : boolean;
  signal type_cast_163_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_988_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_0 : boolean;
  signal WPIPE_Block0_start_988_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 : boolean;
  signal type_cast_610_inst_ack_0 : boolean;
  signal type_cast_610_inst_req_0 : boolean;
  signal type_cast_176_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1051_inst_ack_0 : boolean;
  signal type_cast_176_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_1 : boolean;
  signal type_cast_176_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 : boolean;
  signal type_cast_188_inst_req_0 : boolean;
  signal type_cast_188_inst_ack_0 : boolean;
  signal type_cast_188_inst_req_1 : boolean;
  signal WPIPE_Block0_start_988_inst_ack_1 : boolean;
  signal type_cast_188_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1014_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 : boolean;
  signal type_cast_201_inst_req_0 : boolean;
  signal type_cast_201_inst_ack_0 : boolean;
  signal type_cast_201_inst_req_1 : boolean;
  signal type_cast_201_inst_ack_1 : boolean;
  signal type_cast_210_inst_req_0 : boolean;
  signal type_cast_210_inst_ack_0 : boolean;
  signal type_cast_210_inst_req_1 : boolean;
  signal type_cast_210_inst_ack_1 : boolean;
  signal type_cast_556_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1058_inst_req_1 : boolean;
  signal type_cast_556_inst_req_1 : boolean;
  signal type_cast_214_inst_req_0 : boolean;
  signal type_cast_214_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 : boolean;
  signal type_cast_214_inst_req_1 : boolean;
  signal type_cast_214_inst_ack_1 : boolean;
  signal if_stmt_632_branch_ack_0 : boolean;
  signal type_cast_218_inst_req_0 : boolean;
  signal type_cast_218_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_0 : boolean;
  signal type_cast_218_inst_req_1 : boolean;
  signal type_cast_218_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_997_inst_ack_0 : boolean;
  signal type_cast_556_inst_ack_0 : boolean;
  signal type_cast_556_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1017_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1017_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_ack_1 : boolean;
  signal type_cast_255_inst_req_0 : boolean;
  signal type_cast_255_inst_ack_0 : boolean;
  signal type_cast_255_inst_req_1 : boolean;
  signal type_cast_255_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_req_1 : boolean;
  signal type_cast_259_inst_req_0 : boolean;
  signal type_cast_259_inst_ack_0 : boolean;
  signal type_cast_259_inst_req_1 : boolean;
  signal type_cast_259_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1058_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_ack_0 : boolean;
  signal type_cast_263_inst_req_0 : boolean;
  signal type_cast_263_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1058_inst_req_0 : boolean;
  signal type_cast_263_inst_req_1 : boolean;
  signal type_cast_263_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_req_0 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal type_cast_267_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1051_inst_req_1 : boolean;
  signal type_cast_267_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_req_1 : boolean;
  signal WPIPE_Block0_start_988_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_ack_1 : boolean;
  signal type_cast_709_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1029_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_982_inst_req_1 : boolean;
  signal type_cast_289_inst_req_0 : boolean;
  signal type_cast_289_inst_ack_0 : boolean;
  signal type_cast_289_inst_req_1 : boolean;
  signal type_cast_289_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_ack_0 : boolean;
  signal type_cast_709_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_ack_1 : boolean;
  signal type_cast_302_inst_req_0 : boolean;
  signal type_cast_302_inst_ack_0 : boolean;
  signal type_cast_302_inst_req_1 : boolean;
  signal type_cast_302_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1029_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_ack_1 : boolean;
  signal type_cast_709_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1064_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_ack_1 : boolean;
  signal type_cast_592_inst_ack_1 : boolean;
  signal type_cast_592_inst_req_1 : boolean;
  signal type_cast_314_inst_req_0 : boolean;
  signal type_cast_314_inst_ack_0 : boolean;
  signal type_cast_314_inst_req_1 : boolean;
  signal type_cast_314_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_ack_1 : boolean;
  signal type_cast_327_inst_req_0 : boolean;
  signal type_cast_327_inst_ack_0 : boolean;
  signal type_cast_327_inst_req_1 : boolean;
  signal type_cast_327_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1017_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1017_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1051_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_ack_1 : boolean;
  signal type_cast_352_inst_req_0 : boolean;
  signal type_cast_352_inst_ack_0 : boolean;
  signal type_cast_352_inst_req_1 : boolean;
  signal type_cast_352_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_991_inst_req_1 : boolean;
  signal type_cast_1431_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1076_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_ack_1 : boolean;
  signal type_cast_364_inst_req_0 : boolean;
  signal type_cast_364_inst_ack_0 : boolean;
  signal type_cast_364_inst_req_1 : boolean;
  signal type_cast_364_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_991_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_ack_1 : boolean;
  signal type_cast_377_inst_req_0 : boolean;
  signal type_cast_377_inst_ack_0 : boolean;
  signal type_cast_377_inst_req_1 : boolean;
  signal type_cast_377_inst_ack_1 : boolean;
  signal type_cast_1401_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1020_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1020_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1020_inst_req_1 : boolean;
  signal type_cast_389_inst_req_0 : boolean;
  signal type_cast_389_inst_ack_0 : boolean;
  signal type_cast_389_inst_req_1 : boolean;
  signal type_cast_389_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_req_1 : boolean;
  signal type_cast_1401_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1020_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_976_inst_req_0 : boolean;
  signal type_cast_402_inst_req_0 : boolean;
  signal type_cast_402_inst_ack_0 : boolean;
  signal type_cast_402_inst_req_1 : boolean;
  signal type_cast_402_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_997_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1032_inst_req_0 : boolean;
  signal WPIPE_Block0_start_994_inst_req_0 : boolean;
  signal if_stmt_416_branch_req_0 : boolean;
  signal if_stmt_416_branch_ack_1 : boolean;
  signal if_stmt_416_branch_ack_0 : boolean;
  signal if_stmt_431_branch_req_0 : boolean;
  signal if_stmt_431_branch_ack_1 : boolean;
  signal if_stmt_431_branch_ack_0 : boolean;
  signal type_cast_452_inst_req_0 : boolean;
  signal type_cast_452_inst_ack_0 : boolean;
  signal type_cast_452_inst_req_1 : boolean;
  signal type_cast_452_inst_ack_1 : boolean;
  signal array_obj_ref_481_index_offset_req_0 : boolean;
  signal array_obj_ref_481_index_offset_ack_0 : boolean;
  signal array_obj_ref_481_index_offset_req_1 : boolean;
  signal array_obj_ref_481_index_offset_ack_1 : boolean;
  signal addr_of_482_final_reg_req_0 : boolean;
  signal addr_of_482_final_reg_ack_0 : boolean;
  signal addr_of_482_final_reg_req_1 : boolean;
  signal addr_of_482_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_ack_1 : boolean;
  signal type_cast_489_inst_req_0 : boolean;
  signal type_cast_489_inst_ack_0 : boolean;
  signal type_cast_489_inst_req_1 : boolean;
  signal type_cast_489_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1014_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_ack_1 : boolean;
  signal type_cast_502_inst_req_0 : boolean;
  signal type_cast_502_inst_ack_0 : boolean;
  signal type_cast_502_inst_req_1 : boolean;
  signal type_cast_502_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_ack_1 : boolean;
  signal type_cast_520_inst_req_0 : boolean;
  signal type_cast_520_inst_ack_0 : boolean;
  signal type_cast_520_inst_req_1 : boolean;
  signal type_cast_520_inst_ack_1 : boolean;
  signal type_cast_745_inst_req_0 : boolean;
  signal type_cast_745_inst_ack_0 : boolean;
  signal type_cast_745_inst_req_1 : boolean;
  signal type_cast_745_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1082_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1076_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 : boolean;
  signal type_cast_1431_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_req_1 : boolean;
  signal type_cast_763_inst_req_0 : boolean;
  signal type_cast_1049_inst_ack_1 : boolean;
  signal type_cast_763_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1 : boolean;
  signal type_cast_763_inst_req_1 : boolean;
  signal type_cast_1049_inst_req_1 : boolean;
  signal type_cast_763_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1082_inst_req_0 : boolean;
  signal WPIPE_Block0_start_985_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1061_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1061_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1076_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_985_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1008_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1070_inst_ack_1 : boolean;
  signal type_cast_781_inst_req_0 : boolean;
  signal type_cast_1049_inst_ack_0 : boolean;
  signal type_cast_781_inst_ack_0 : boolean;
  signal type_cast_781_inst_req_1 : boolean;
  signal type_cast_1049_inst_req_0 : boolean;
  signal type_cast_781_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 : boolean;
  signal type_cast_1431_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1008_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1070_inst_req_1 : boolean;
  signal type_cast_799_inst_req_0 : boolean;
  signal type_cast_799_inst_ack_0 : boolean;
  signal type_cast_799_inst_req_1 : boolean;
  signal type_cast_799_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_985_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1008_inst_ack_0 : boolean;
  signal type_cast_817_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1038_inst_ack_1 : boolean;
  signal type_cast_817_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1067_inst_ack_1 : boolean;
  signal type_cast_817_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1038_inst_req_1 : boolean;
  signal type_cast_817_inst_ack_1 : boolean;
  signal type_cast_1056_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1008_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1038_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1038_inst_req_0 : boolean;
  signal ptr_deref_825_store_0_req_0 : boolean;
  signal ptr_deref_825_store_0_ack_0 : boolean;
  signal ptr_deref_825_store_0_req_1 : boolean;
  signal ptr_deref_825_store_0_ack_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1073_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1067_inst_req_1 : boolean;
  signal WPIPE_Block0_start_979_inst_ack_1 : boolean;
  signal if_stmt_839_branch_req_0 : boolean;
  signal WPIPE_Block0_start_1005_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_979_inst_req_1 : boolean;
  signal if_stmt_839_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1026_inst_ack_1 : boolean;
  signal if_stmt_839_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1026_inst_req_1 : boolean;
  signal type_cast_1056_inst_req_1 : boolean;
  signal type_cast_850_inst_req_0 : boolean;
  signal type_cast_850_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1 : boolean;
  signal type_cast_850_inst_req_1 : boolean;
  signal type_cast_850_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1073_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_req_0 : boolean;
  signal type_cast_1371_inst_req_0 : boolean;
  signal array_obj_ref_1362_index_offset_req_1 : boolean;
  signal WPIPE_Block0_start_1005_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1067_inst_ack_0 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal type_cast_854_inst_req_1 : boolean;
  signal type_cast_854_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1085_inst_req_1 : boolean;
  signal type_cast_1056_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1067_inst_req_0 : boolean;
  signal type_cast_858_inst_req_0 : boolean;
  signal type_cast_858_inst_ack_0 : boolean;
  signal type_cast_858_inst_req_1 : boolean;
  signal type_cast_858_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1073_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_979_inst_ack_0 : boolean;
  signal if_stmt_876_branch_req_0 : boolean;
  signal WPIPE_Block0_start_979_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1026_inst_ack_0 : boolean;
  signal if_stmt_876_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1026_inst_req_0 : boolean;
  signal if_stmt_876_branch_ack_0 : boolean;
  signal WPIPE_Block2_start_1082_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_994_inst_ack_1 : boolean;
  signal type_cast_903_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1035_inst_ack_1 : boolean;
  signal type_cast_903_inst_ack_0 : boolean;
  signal type_cast_903_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1035_inst_req_1 : boolean;
  signal type_cast_903_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1073_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0 : boolean;
  signal type_cast_1371_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1070_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1064_inst_ack_0 : boolean;
  signal type_cast_1056_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1005_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1064_inst_req_0 : boolean;
  signal array_obj_ref_1362_index_offset_ack_1 : boolean;
  signal WPIPE_Block2_start_1079_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1005_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1 : boolean;
  signal array_obj_ref_932_index_offset_req_0 : boolean;
  signal array_obj_ref_932_index_offset_ack_0 : boolean;
  signal WPIPE_Block0_start_985_inst_req_0 : boolean;
  signal array_obj_ref_932_index_offset_req_1 : boolean;
  signal array_obj_ref_932_index_offset_ack_1 : boolean;
  signal WPIPE_Block1_start_1035_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1035_inst_req_0 : boolean;
  signal addr_of_933_final_reg_req_0 : boolean;
  signal addr_of_933_final_reg_ack_0 : boolean;
  signal addr_of_933_final_reg_req_1 : boolean;
  signal addr_of_933_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1079_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1023_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_994_inst_req_1 : boolean;
  signal ptr_deref_936_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1001_inst_ack_1 : boolean;
  signal ptr_deref_936_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1023_inst_req_1 : boolean;
  signal ptr_deref_936_store_0_req_1 : boolean;
  signal WPIPE_Block0_start_1001_inst_req_1 : boolean;
  signal ptr_deref_936_store_0_ack_1 : boolean;
  signal WPIPE_Block2_start_1076_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1082_inst_req_1 : boolean;
  signal if_stmt_951_branch_req_0 : boolean;
  signal WPIPE_Block2_start_1070_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1001_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_1 : boolean;
  signal if_stmt_951_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1023_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_976_inst_req_1 : boolean;
  signal if_stmt_951_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_994_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1023_inst_req_0 : boolean;
  signal type_cast_1371_inst_req_1 : boolean;
  signal call_stmt_962_call_req_0 : boolean;
  signal WPIPE_Block1_start_1032_inst_ack_1 : boolean;
  signal call_stmt_962_call_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1 : boolean;
  signal call_stmt_962_call_req_1 : boolean;
  signal WPIPE_Block1_start_1032_inst_req_1 : boolean;
  signal call_stmt_962_call_ack_1 : boolean;
  signal type_cast_1401_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1001_inst_req_0 : boolean;
  signal type_cast_967_inst_req_0 : boolean;
  signal type_cast_967_inst_ack_0 : boolean;
  signal type_cast_967_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1032_inst_ack_0 : boolean;
  signal type_cast_967_inst_ack_1 : boolean;
  signal type_cast_1381_inst_req_0 : boolean;
  signal array_obj_ref_1362_index_offset_req_0 : boolean;
  signal WPIPE_Block0_start_970_inst_req_0 : boolean;
  signal WPIPE_Block0_start_970_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_970_inst_req_1 : boolean;
  signal WPIPE_Block0_start_970_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1088_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1088_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1088_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1091_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1091_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1091_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1094_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1094_inst_ack_1 : boolean;
  signal type_cast_1105_inst_req_0 : boolean;
  signal ptr_deref_1367_load_0_ack_1 : boolean;
  signal type_cast_1105_inst_ack_0 : boolean;
  signal type_cast_1441_inst_ack_1 : boolean;
  signal type_cast_1105_inst_req_1 : boolean;
  signal ptr_deref_1367_load_0_req_1 : boolean;
  signal type_cast_1105_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1107_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1107_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1107_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1107_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1446_inst_ack_1 : boolean;
  signal type_cast_1391_inst_ack_1 : boolean;
  signal type_cast_1391_inst_req_1 : boolean;
  signal type_cast_1441_inst_req_1 : boolean;
  signal type_cast_1112_inst_req_0 : boolean;
  signal type_cast_1112_inst_ack_0 : boolean;
  signal type_cast_1112_inst_req_1 : boolean;
  signal type_cast_1112_inst_ack_1 : boolean;
  signal type_cast_1421_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1114_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1114_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1114_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1114_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1446_inst_req_1 : boolean;
  signal type_cast_1391_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1117_inst_req_0 : boolean;
  signal ptr_deref_1367_load_0_ack_0 : boolean;
  signal WPIPE_Block2_start_1117_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1117_inst_req_1 : boolean;
  signal ptr_deref_1367_load_0_req_0 : boolean;
  signal WPIPE_Block2_start_1117_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_req_0 : boolean;
  signal type_cast_1391_inst_req_0 : boolean;
  signal type_cast_1421_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1120_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1120_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1120_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1120_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1446_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1123_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1123_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1123_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1123_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1446_inst_req_0 : boolean;
  signal type_cast_1333_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1126_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1126_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1126_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1126_inst_ack_1 : boolean;
  signal type_cast_1333_inst_req_1 : boolean;
  signal type_cast_1421_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1129_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1129_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1129_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1129_inst_ack_1 : boolean;
  signal type_cast_1421_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1132_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1132_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1132_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1132_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1135_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1135_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1135_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1135_inst_ack_1 : boolean;
  signal type_cast_1333_inst_ack_0 : boolean;
  signal type_cast_1333_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1138_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1138_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1138_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1138_inst_ack_1 : boolean;
  signal type_cast_1381_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1141_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1141_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1141_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1141_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1144_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1144_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1144_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1144_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1443_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1147_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1147_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1147_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1147_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1443_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1150_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1150_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1150_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1150_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1443_inst_ack_0 : boolean;
  signal if_stmt_1306_branch_ack_0 : boolean;
  signal type_cast_1161_inst_req_0 : boolean;
  signal type_cast_1161_inst_ack_0 : boolean;
  signal type_cast_1441_inst_ack_0 : boolean;
  signal type_cast_1161_inst_req_1 : boolean;
  signal type_cast_1161_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_0 : boolean;
  signal type_cast_1381_inst_req_1 : boolean;
  signal if_stmt_1306_branch_ack_1 : boolean;
  signal type_cast_1411_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1163_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1163_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1163_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1163_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1443_inst_req_0 : boolean;
  signal if_stmt_1306_branch_req_0 : boolean;
  signal type_cast_1441_inst_req_0 : boolean;
  signal type_cast_1168_inst_req_0 : boolean;
  signal addr_of_1363_final_reg_ack_1 : boolean;
  signal type_cast_1168_inst_ack_0 : boolean;
  signal type_cast_1168_inst_req_1 : boolean;
  signal addr_of_1363_final_reg_req_1 : boolean;
  signal type_cast_1168_inst_ack_1 : boolean;
  signal type_cast_1381_inst_ack_0 : boolean;
  signal type_cast_1411_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1170_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1170_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1170_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1170_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1173_inst_req_0 : boolean;
  signal addr_of_1363_final_reg_ack_0 : boolean;
  signal WPIPE_Block3_start_1173_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1173_inst_req_1 : boolean;
  signal addr_of_1363_final_reg_req_0 : boolean;
  signal WPIPE_Block3_start_1173_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1176_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1176_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1176_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1176_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0 : boolean;
  signal type_cast_1411_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1179_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1179_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1179_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1179_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_req_0 : boolean;
  signal type_cast_1411_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1183_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1183_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1183_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1183_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1186_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1186_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1186_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1186_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1189_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1189_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1189_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1189_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1192_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1192_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1192_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1192_inst_ack_1 : boolean;
  signal call_stmt_1196_call_req_0 : boolean;
  signal call_stmt_1196_call_ack_0 : boolean;
  signal call_stmt_1196_call_req_1 : boolean;
  signal call_stmt_1196_call_ack_1 : boolean;
  signal type_cast_1200_inst_req_0 : boolean;
  signal type_cast_1200_inst_ack_0 : boolean;
  signal type_cast_1200_inst_req_1 : boolean;
  signal type_cast_1200_inst_ack_1 : boolean;
  signal type_cast_1209_inst_req_0 : boolean;
  signal type_cast_1209_inst_ack_0 : boolean;
  signal type_cast_1209_inst_req_1 : boolean;
  signal type_cast_1209_inst_ack_1 : boolean;
  signal type_cast_1219_inst_req_0 : boolean;
  signal type_cast_1219_inst_ack_0 : boolean;
  signal type_cast_1219_inst_req_1 : boolean;
  signal type_cast_1219_inst_ack_1 : boolean;
  signal type_cast_1229_inst_req_0 : boolean;
  signal type_cast_1229_inst_ack_0 : boolean;
  signal type_cast_1229_inst_req_1 : boolean;
  signal type_cast_1229_inst_ack_1 : boolean;
  signal type_cast_1239_inst_req_0 : boolean;
  signal type_cast_1239_inst_ack_0 : boolean;
  signal type_cast_1239_inst_req_1 : boolean;
  signal type_cast_1239_inst_ack_1 : boolean;
  signal type_cast_1249_inst_req_0 : boolean;
  signal type_cast_1249_inst_ack_0 : boolean;
  signal type_cast_1249_inst_req_1 : boolean;
  signal type_cast_1249_inst_ack_1 : boolean;
  signal type_cast_1259_inst_req_0 : boolean;
  signal type_cast_1259_inst_ack_0 : boolean;
  signal type_cast_1259_inst_req_1 : boolean;
  signal type_cast_1259_inst_ack_1 : boolean;
  signal type_cast_1269_inst_req_0 : boolean;
  signal type_cast_1269_inst_ack_0 : boolean;
  signal type_cast_1269_inst_req_1 : boolean;
  signal type_cast_1269_inst_ack_1 : boolean;
  signal type_cast_1279_inst_req_0 : boolean;
  signal type_cast_1279_inst_ack_0 : boolean;
  signal type_cast_1279_inst_req_1 : boolean;
  signal type_cast_1279_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1 : boolean;
  signal if_stmt_1478_branch_req_0 : boolean;
  signal if_stmt_1478_branch_ack_1 : boolean;
  signal if_stmt_1478_branch_ack_0 : boolean;
  signal phi_stmt_469_req_0 : boolean;
  signal type_cast_475_inst_req_0 : boolean;
  signal type_cast_475_inst_ack_0 : boolean;
  signal type_cast_475_inst_req_1 : boolean;
  signal type_cast_475_inst_ack_1 : boolean;
  signal phi_stmt_469_req_1 : boolean;
  signal phi_stmt_469_ack_0 : boolean;
  signal phi_stmt_676_req_1 : boolean;
  signal type_cast_679_inst_req_0 : boolean;
  signal type_cast_679_inst_ack_0 : boolean;
  signal type_cast_679_inst_req_1 : boolean;
  signal type_cast_679_inst_ack_1 : boolean;
  signal phi_stmt_676_req_0 : boolean;
  signal phi_stmt_676_ack_0 : boolean;
  signal phi_stmt_920_req_1 : boolean;
  signal type_cast_923_inst_req_0 : boolean;
  signal type_cast_923_inst_ack_0 : boolean;
  signal type_cast_923_inst_req_1 : boolean;
  signal type_cast_923_inst_ack_1 : boolean;
  signal phi_stmt_920_req_0 : boolean;
  signal phi_stmt_920_ack_0 : boolean;
  signal phi_stmt_1350_req_0 : boolean;
  signal type_cast_1356_inst_req_0 : boolean;
  signal type_cast_1356_inst_ack_0 : boolean;
  signal type_cast_1356_inst_req_1 : boolean;
  signal type_cast_1356_inst_ack_1 : boolean;
  signal phi_stmt_1350_req_1 : boolean;
  signal phi_stmt_1350_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(496 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(496);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/cr
      -- 
    rr_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_51_inst_req_1); -- 
    cr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_63_inst_req_1); -- 
    cr_238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_76_inst_req_1); -- 
    cr_266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_88_inst_req_1); -- 
    cr_294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_101_inst_req_1); -- 
    cr_322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_113_inst_req_1); -- 
    cr_350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_126_inst_req_1); -- 
    cr_756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_339_inst_req_1); -- 
    cr_378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_138_inst_req_1); -- 
    cr_406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_151_inst_req_1); -- 
    cr_434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_163_inst_req_1); -- 
    cr_462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_176_inst_req_1); -- 
    cr_490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_188_inst_req_1); -- 
    cr_518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_201_inst_req_1); -- 
    cr_532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_210_inst_req_1); -- 
    cr_546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_214_inst_req_1); -- 
    cr_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_218_inst_req_1); -- 
    cr_574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_255_inst_req_1); -- 
    cr_588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_259_inst_req_1); -- 
    cr_602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_263_inst_req_1); -- 
    cr_616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_267_inst_req_1); -- 
    cr_644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_289_inst_req_1); -- 
    cr_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_302_inst_req_1); -- 
    cr_700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_314_inst_req_1); -- 
    cr_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_327_inst_req_1); -- 
    cr_784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_352_inst_req_1); -- 
    cr_812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_364_inst_req_1); -- 
    cr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_377_inst_req_1); -- 
    cr_868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_389_inst_req_1); -- 
    cr_896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_402_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/rr
      -- 
    ca_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/ra
      -- 
    ra_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/ca
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_update_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/cr
      -- 
    ra_164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/rr
      -- 
    ca_169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_51_inst_req_0); -- 
    rr_191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/ra
      -- 
    ra_178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/ca
      -- 
    ca_183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_update_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/cr
      -- 
    ra_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/rr
      -- 
    ca_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_63_inst_req_0); -- 
    rr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/ra
      -- 
    ra_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/ca
      -- 
    ca_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_update_start_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/cr
      -- 
    ra_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/rr
      -- 
    ca_225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_76_inst_req_0); -- 
    rr_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/ra
      -- 
    ra_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/ca
      -- 
    ca_239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_update_start_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/cr
      -- 
    ra_248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/rr
      -- 
    ca_253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_88_inst_req_0); -- 
    rr_275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/ra
      -- 
    ra_262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/ca
      -- 
    ca_267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_update_start_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/cr
      -- 
    ra_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/rr
      -- 
    ca_281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_101_inst_req_0); -- 
    rr_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/ra
      -- 
    ra_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/ca
      -- 
    ca_295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_update_start_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/cr
      -- 
    ra_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/rr
      -- 
    ca_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_113_inst_req_0); -- 
    rr_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/ra
      -- 
    ra_318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/ca
      -- 
    ca_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_update_start_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/cr
      -- 
    ra_332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/$entry
      -- 
    ca_337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_126_inst_req_0); -- 
    rr_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/ra
      -- 
    ra_346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/ca
      -- 
    ca_351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_update_start_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/$exit
      -- 
    ra_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/rr
      -- 
    ca_365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_138_inst_req_0); -- 
    rr_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/ra
      -- 
    ra_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/ca
      -- 
    ca_379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_update_start_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/cr
      -- 
    ra_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/rr
      -- 
    ca_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_0); -- 
    rr_401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_151_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/ra
      -- 
    ra_402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/ca
      -- 
    ca_407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_update_start_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/cr
      -- 
    ra_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/rr
      -- 
    ca_421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_163_inst_req_0); -- 
    rr_443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/ra
      -- 
    ra_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/ca
      -- 
    ca_435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_update_start_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/cr
      -- 
    ra_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/rr
      -- 
    ca_449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_0); -- 
    rr_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_176_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/ra
      -- 
    ra_458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/ca
      -- 
    ca_463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_update_start_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/cr
      -- 
    ra_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/rr
      -- 
    ca_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_188_inst_req_0); -- 
    rr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/ra
      -- 
    ra_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/ca
      -- 
    ca_491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_update_start_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/cr
      -- 
    ra_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/rr
      -- 
    ca_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_201_inst_req_0); -- 
    rr_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_285_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/ra
      -- 
    ra_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/ca
      -- 
    ca_519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/rr
      -- 
    rr_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_210_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/ra
      -- 
    ra_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_0, ack => convTranspose_CP_39_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/ca
      -- 
    ca_533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_1, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/rr
      -- 
    rr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => type_cast_214_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/ra
      -- 
    ra_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/ca
      -- 
    ca_547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/rr
      -- 
    rr_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => type_cast_218_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/ra
      -- 
    ra_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_0, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/ca
      -- 
    ca_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_1, ack => convTranspose_CP_39_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/rr
      -- 
    rr_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_255_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/ra
      -- 
    ra_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/ca
      -- 
    ca_575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/rr
      -- 
    rr_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => type_cast_259_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/ra
      -- 
    ra_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_259_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/ca
      -- 
    ca_589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_259_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	48 
    -- CP-element group 72: 	44 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/rr
      -- 
    rr_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => type_cast_263_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(48) & convTranspose_CP_39_elements(44);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/ra
      -- 
    ra_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/ca
      -- 
    ca_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	56 
    -- CP-element group 75: 	52 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/rr
      -- 
    rr_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(75), ack => type_cast_267_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(56) & convTranspose_CP_39_elements(52);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/ra
      -- 
    ra_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_0, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/ca
      -- 
    ca_617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_1, ack => convTranspose_CP_39_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_update_start_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/cr
      -- 
    ra_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_285_inst_ack_0, ack => convTranspose_CP_39_elements(78)); -- 
    cr_630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_285_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/rr
      -- 
    ca_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_285_inst_ack_1, ack => convTranspose_CP_39_elements(79)); -- 
    rr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => type_cast_289_inst_req_0); -- 
    rr_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => RPIPE_ConvTranspose_input_pipe_298_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/ra
      -- 
    ra_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_289_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/ca
      -- 
    ca_645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_289_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_update_start_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/cr
      -- 
    ra_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_298_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    cr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_298_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/rr
      -- 
    ca_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_298_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    rr_667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => type_cast_302_inst_req_0); -- 
    rr_681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => RPIPE_ConvTranspose_input_pipe_310_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/ra
      -- 
    ra_668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/ca
      -- 
    ca_673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_update_start_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/cr
      -- 
    ra_682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_310_inst_ack_0, ack => convTranspose_CP_39_elements(86)); -- 
    cr_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_310_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/rr
      -- 
    ca_687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_310_inst_ack_1, ack => convTranspose_CP_39_elements(87)); -- 
    rr_695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => type_cast_314_inst_req_0); -- 
    rr_709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => RPIPE_ConvTranspose_input_pipe_323_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/ra
      -- 
    ra_696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_314_inst_ack_0, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/ca
      -- 
    ca_701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_314_inst_ack_1, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_update_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/cr
      -- 
    ra_710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_323_inst_ack_0, ack => convTranspose_CP_39_elements(90)); -- 
    cr_714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_323_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/rr
      -- 
    ca_715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_323_inst_ack_1, ack => convTranspose_CP_39_elements(91)); -- 
    rr_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => type_cast_327_inst_req_0); -- 
    rr_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_335_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/ra
      -- 
    ra_724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_327_inst_ack_0, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/ca
      -- 
    ca_729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_327_inst_ack_1, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_update_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/cr
      -- 
    ra_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_335_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    cr_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => RPIPE_ConvTranspose_input_pipe_335_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_sample_start_
      -- 
    ca_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_335_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    rr_751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => type_cast_339_inst_req_0); -- 
    rr_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => RPIPE_ConvTranspose_input_pipe_348_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_sample_completed_
      -- 
    ra_752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_update_completed_
      -- 
    ca_757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_update_start_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/cr
      -- 
    ra_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_348_inst_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    cr_770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => RPIPE_ConvTranspose_input_pipe_348_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/rr
      -- 
    ca_771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_348_inst_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    rr_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => type_cast_352_inst_req_0); -- 
    rr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => RPIPE_ConvTranspose_input_pipe_360_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/ra
      -- 
    ra_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/ca
      -- 
    ca_785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_update_start_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/cr
      -- 
    ra_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_360_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    cr_798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(102), ack => RPIPE_ConvTranspose_input_pipe_360_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/rr
      -- 
    ca_799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_360_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    rr_807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => type_cast_364_inst_req_0); -- 
    rr_821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => RPIPE_ConvTranspose_input_pipe_373_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/ra
      -- 
    ra_808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_364_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/ca
      -- 
    ca_813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_364_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_update_start_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/cr
      -- 
    ra_822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_373_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    cr_826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(106), ack => RPIPE_ConvTranspose_input_pipe_373_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/rr
      -- 
    ca_827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_373_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    rr_835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_377_inst_req_0); -- 
    rr_849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => RPIPE_ConvTranspose_input_pipe_385_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/ra
      -- 
    ra_836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_377_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/ca
      -- 
    ca_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_377_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_update_start_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/cr
      -- 
    ra_850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_385_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    cr_854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => RPIPE_ConvTranspose_input_pipe_385_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/rr
      -- 
    ca_855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_385_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    rr_863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => type_cast_389_inst_req_0); -- 
    rr_877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => RPIPE_ConvTranspose_input_pipe_398_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/ra
      -- 
    ra_864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_389_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/ca
      -- 
    ca_869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_389_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_update_start_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/cr
      -- 
    ra_878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_398_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    cr_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(114), ack => RPIPE_ConvTranspose_input_pipe_398_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/rr
      -- 
    ca_883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_398_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    rr_891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(115), ack => type_cast_402_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/ra
      -- 
    ra_892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/ca
      -- 
    ca_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415__exit__
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416__entry__
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_32/R_cmp513_417_place
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_else_link/$entry
      -- 
    branch_req_905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(118), ack => if_stmt_416_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(59) & convTranspose_CP_39_elements(62) & convTranspose_CP_39_elements(65) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(77) & convTranspose_CP_39_elements(81) & convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(89) & convTranspose_CP_39_elements(93) & convTranspose_CP_39_elements(97) & convTranspose_CP_39_elements(101) & convTranspose_CP_39_elements(105) & convTranspose_CP_39_elements(109) & convTranspose_CP_39_elements(113) & convTranspose_CP_39_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437__exit__
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466__entry__
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_416_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_416_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph515
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_update_start_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph515_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph515_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/dummy
      -- 
    if_choice_transition_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_416_branch_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    rr_949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_452_inst_req_0); -- 
    cr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_452_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	469 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_416_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_416_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_416_branch_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	469 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638__exit__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673__entry__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_update_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_431_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_431_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph511
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/dummy
      -- 
    if_choice_transition_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_431_branch_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    cr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_659_inst_req_1); -- 
    rr_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_659_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	469 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	482 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_431_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_431_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_431_branch_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/ra
      -- 
    ra_950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_0, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	470 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466__exit__
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$entry
      -- 
    ca_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_1, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	475 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/ack
      -- 
    ack_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_481_index_offset_ack_0, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	475 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/req
      -- 
    ack_989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_481_index_offset_ack_1, ack => convTranspose_CP_39_elements(126)); -- 
    req_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => addr_of_482_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/ack
      -- 
    ack_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_482_final_reg_ack_0, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	475 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/ack
      -- 
    ack_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_482_final_reg_ack_1, ack => convTranspose_CP_39_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	475 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_update_start_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/cr
      -- 
    ra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_485_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    cr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_485_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/rr
      -- 
    ca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_485_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    rr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => type_cast_489_inst_req_0); -- 
    rr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => RPIPE_ConvTranspose_input_pipe_498_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/ra
      -- 
    ra_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_489_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	475 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/ca
      -- 
    ca_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_489_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_update_start_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/cr
      -- 
    ra_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_498_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_498_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/rr
      -- 
    ca_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_498_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_502_inst_req_0); -- 
    rr_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_516_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/ra
      -- 
    ra_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_0, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	475 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/ca
      -- 
    ca_1060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_update_start_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/cr
      -- 
    ra_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_516_inst_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    cr_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => RPIPE_ConvTranspose_input_pipe_516_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_sample_start_
      -- 
    ca_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_516_inst_ack_1, ack => convTranspose_CP_39_elements(138)); -- 
    rr_1082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => type_cast_520_inst_req_0); -- 
    rr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/ra
      -- 
    ra_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_0, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	475 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/ca
      -- 
    ca_1088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_1, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_update_start_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_sample_completed_
      -- 
    ra_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    cr_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_sample_start_
      -- 
    ca_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    rr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => type_cast_538_inst_req_0); -- 
    rr_1124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => RPIPE_ConvTranspose_input_pipe_552_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_sample_completed_
      -- 
    ra_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	475 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_update_completed_
      -- 
    ca_1116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_update_start_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_sample_completed_
      -- 
    ra_1125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_552_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    cr_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_552_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_update_completed_
      -- 
    ca_1130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_552_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    rr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => type_cast_556_inst_req_0); -- 
    rr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => RPIPE_ConvTranspose_input_pipe_570_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_sample_completed_
      -- 
    ra_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	475 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_update_completed_
      -- 
    ca_1144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_update_start_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_sample_completed_
      -- 
    ra_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_570_inst_ack_0, ack => convTranspose_CP_39_elements(149)); -- 
    cr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_570_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_update_completed_
      -- 
    ca_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_570_inst_ack_1, ack => convTranspose_CP_39_elements(150)); -- 
    rr_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => type_cast_574_inst_req_0); -- 
    rr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => RPIPE_ConvTranspose_input_pipe_588_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_sample_completed_
      -- 
    ra_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_0, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	475 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_update_completed_
      -- 
    ca_1172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_1, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_update_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_sample_completed_
      -- 
    ra_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_588_inst_ack_0, ack => convTranspose_CP_39_elements(153)); -- 
    cr_1185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_588_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	157 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_sample_start_
      -- 
    ca_1186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_588_inst_ack_1, ack => convTranspose_CP_39_elements(154)); -- 
    rr_1194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => type_cast_592_inst_req_0); -- 
    rr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_606_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_sample_completed_
      -- 
    ra_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_0, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	475 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/ca
      -- 
    ca_1200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_1, ack => convTranspose_CP_39_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_update_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_sample_completed_
      -- 
    ra_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_606_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_606_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_update_completed_
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_606_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    rr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(158), ack => type_cast_610_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_sample_completed_
      -- 
    ra_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	475 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_update_completed_
      -- 
    ca_1228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/$entry
      -- 
    rr_1266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => ptr_deref_618_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(160) & convTranspose_CP_39_elements(128) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(136) & convTranspose_CP_39_elements(140) & convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(152) & convTranspose_CP_39_elements(156);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/$exit
      -- 
    ra_1267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_618_store_0_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	475 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_update_completed_
      -- 
    ca_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_618_store_0_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631__exit__
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632__entry__
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/R_exitcond3_633_place
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/$exit
      -- 
    branch_req_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => if_stmt_632_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	469 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422__exit__
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_632_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_632_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_632_branch_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	471 
    -- CP-element group 166: 	472 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_632_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_632_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_632_branch_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    rr_3511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_475_inst_req_0); -- 
    cr_3516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_475_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_sample_completed_
      -- 
    ra_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_0, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	476 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673__exit__
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$entry
      -- 
    ca_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_1, ack => convTranspose_CP_39_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	481 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_sample_complete
      -- 
    ack_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_index_offset_ack_0, ack => convTranspose_CP_39_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	481 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/req
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/sum_rename_ack
      -- 
    ack_1348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_index_offset_ack_1, ack => convTranspose_CP_39_elements(170)); -- 
    req_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => addr_of_689_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/ack
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/$exit
      -- 
    ack_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_689_final_reg_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	481 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/root_register_ack
      -- 
    ack_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_689_final_reg_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	481 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_update_start_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_sample_completed_
      -- 
    ra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_692_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    cr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_692_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/ca
      -- 
    ca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_692_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    rr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => type_cast_696_inst_req_0); -- 
    rr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_sample_completed_
      -- 
    ra_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_696_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	481 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_update_completed_
      -- 
    ca_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_696_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_update_start_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/$entry
      -- 
    ra_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/rr
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_0); -- 
    rr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => type_cast_709_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_sample_completed_
      -- 
    ra_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_0, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	481 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/ca
      -- 
    ca_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_update_start_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_sample_completed_
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/$entry
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_727_inst_req_0); -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_sample_completed_
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	481 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/ca
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_update_start_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/cr
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/rr
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => type_cast_745_inst_req_0); -- 
    rr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/ra
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	481 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/ca
      -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_update_start_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/cr
      -- 
    ra_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/rr
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_763_inst_req_0); -- 
    rr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/ra
      -- 
    ra_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	481 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/ca
      -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_update_start_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/cr
      -- 
    ra_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    cr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(193), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/rr
      -- 
    ca_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_1, ack => convTranspose_CP_39_elements(194)); -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_781_inst_req_0); -- 
    rr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/ra
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	481 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/ca
      -- 
    ca_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_update_start_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/cr
      -- 
    ra_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    cr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/rr
      -- 
    ca_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => type_cast_799_inst_req_0); -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => RPIPE_ConvTranspose_input_pipe_813_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/ra
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	481 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/ca
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_update_start_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/cr
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_813_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_813_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/rr
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_813_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_817_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/ra
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	481 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/ca
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	172 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/rr
      -- 
    rr_1625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => ptr_deref_825_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(184) & convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(192) & convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(176) & convTranspose_CP_39_elements(200) & convTranspose_CP_39_elements(204) & convTranspose_CP_39_elements(172);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/ra
      -- 
    ra_1626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_825_store_0_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	481 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/ca
      -- 
    ca_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_825_store_0_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838__exit__
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839__entry__
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_32/R_exitcond2_840_place
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_else_link/$entry
      -- 
    branch_req_1645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => if_stmt_839_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(207) & convTranspose_CP_39_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	482 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845__exit__
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_839_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_839_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_839_branch_ack_1, ack => convTranspose_CP_39_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	477 
    -- CP-element group 210: 	478 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_839_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_839_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_839_branch_ack_0, ack => convTranspose_CP_39_elements(210)); -- 
    rr_3565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_679_inst_req_0); -- 
    cr_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_679_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	482 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/ra
      -- 
    ra_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	482 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/ca
      -- 
    ca_1673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	482 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/ra
      -- 
    ra_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	482 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/ca
      -- 
    ca_1687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	482 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/ra
      -- 
    ra_1696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_858_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	482 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/ca
      -- 
    ca_1701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_858_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875__exit__
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876__entry__
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_32/R_cmp264505_877_place
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_else_link/$entry
      -- 
    branch_req_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => if_stmt_876_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(212) & convTranspose_CP_39_elements(214) & convTranspose_CP_39_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882__exit__
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917__entry__
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_876_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_876_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph507
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_update_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph507_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph507_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/dummy
      -- 
    if_choice_transition_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_876_branch_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    rr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_903_inst_req_0); -- 
    cr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_903_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	489 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_876_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_876_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_876_branch_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/ra
      -- 
    ra_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	483 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917__exit__
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$entry
      -- 
    ca_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	488 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/ack
      -- 
    ack_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_offset_ack_0, ack => convTranspose_CP_39_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	488 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/req
      -- 
    ack_1771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_offset_ack_1, ack => convTranspose_CP_39_elements(223)); -- 
    req_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => addr_of_933_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/ack
      -- 
    ack_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_933_final_reg_ack_0, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	488 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/rr
      -- 
    ack_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_933_final_reg_ack_1, ack => convTranspose_CP_39_elements(225)); -- 
    rr_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => ptr_deref_936_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/ra
      -- 
    ra_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_936_store_0_ack_0, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	488 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/ca
      -- 
    ca_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_936_store_0_ack_1, ack => convTranspose_CP_39_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950__exit__
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951__entry__
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_32/R_exitcond_952_place
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_else_link/$entry
      -- 
    branch_req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => if_stmt_951_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(222) & convTranspose_CP_39_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	489 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957__exit__
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_951_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_951_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_951_branch_ack_1, ack => convTranspose_CP_39_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	484 
    -- CP-element group 230: 	485 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_951_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_951_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_951_branch_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    rr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_923_inst_req_0); -- 
    cr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_923_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	489 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_Sample/cra
      -- 
    cra_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_962_call_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	489 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_Sample/rr
      -- 
    cca_1872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_962_call_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    rr_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => type_cast_967_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_Sample/ra
      -- 
    ra_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	489 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	315 
    -- CP-element group 234: 	316 
    -- CP-element group 234: 	320 
    -- CP-element group 234: 	321 
    -- CP-element group 234: 	331 
    -- CP-element group 234: 	349 
    -- CP-element group 234: 	350 
    -- CP-element group 234: 	354 
    -- CP-element group 234: 	355 
    -- CP-element group 234: 	365 
    -- CP-element group 234: 	367 
    -- CP-element group 234: 	369 
    -- CP-element group 234: 	371 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	263 
    -- CP-element group 234: 	281 
    -- CP-element group 234: 	282 
    -- CP-element group 234: 	286 
    -- CP-element group 234: 	287 
    -- CP-element group 234: 	297 
    -- CP-element group 234:  members (67) 
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968__exit__
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193__entry__
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_update_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_update_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_update_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_update_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_update_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_update_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_Sample/rr
      -- 
    ca_1886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block1_start_1014_inst_req_0); -- 
    cr_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1049_inst_req_1); -- 
    rr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1049_inst_req_0); -- 
    cr_2252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1056_inst_req_1); -- 
    rr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1056_inst_req_0); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block2_start_1070_inst_req_0); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block0_start_970_inst_req_0); -- 
    rr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1105_inst_req_0); -- 
    cr_2448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1105_inst_req_1); -- 
    rr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1112_inst_req_0); -- 
    cr_2476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1112_inst_req_1); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block3_start_1126_inst_req_0); -- 
    rr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1161_inst_req_0); -- 
    cr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1161_inst_req_1); -- 
    rr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1168_inst_req_0); -- 
    cr_2700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => type_cast_1168_inst_req_1); -- 
    rr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_Block0_done_1183_inst_req_0); -- 
    rr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_Block1_done_1186_inst_req_0); -- 
    rr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_Block2_done_1189_inst_req_0); -- 
    rr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => RPIPE_Block3_done_1192_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_update_start_
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_Update/req
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_970_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_970_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_970_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_sample_start_
      -- 
    ack_1903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_970_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_973_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_Update/req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_sample_completed_
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_973_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_973_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_973_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_Sample/req
      -- 
    ack_1917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_973_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_976_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_update_start_
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_Update/req
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_976_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_Sample/req
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_976_Update/ack
      -- 
    ack_1931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_979_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_Update/req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_sample_completed_
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_979_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_979_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_979_update_completed_
      -- 
    ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_979_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_982_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_update_start_
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_Update/req
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_982_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_1958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_982_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_982_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_Sample/$entry
      -- 
    ack_1959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_982_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_985_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_update_start_
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_Update/req
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_Sample/$exit
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_985_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_1972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_985_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_985_update_completed_
      -- 
    ack_1973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_985_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_988_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_Update/req
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_sample_completed_
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_988_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_988_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_988_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_Sample/$entry
      -- 
    ack_1987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_988_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_991_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_Update/req
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_991_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_2000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_991_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_991_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_Sample/req
      -- 
    ack_2001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_991_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_994_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_update_start_
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_Update/req
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_Sample/ack
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_994_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_994_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_994_Update/$exit
      -- 
    ack_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_994_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_997_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_Update/req
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_update_start_
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_sample_completed_
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_997_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_997_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_997_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_Sample/$entry
      -- 
    ack_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_997_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block0_start_1001_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_Update/req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_Sample/$exit
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1001_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block0_start_1001_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1001_Update/$exit
      -- 
    ack_2043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1001_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block0_start_1005_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_Update/req
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_update_start_
      -- CP-element group 257: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_sample_completed_
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1005_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block0_start_1005_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1005_update_completed_
      -- 
    ack_2057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1005_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(258), ack => WPIPE_Block0_start_1008_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_Update/req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_sample_completed_
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1008_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block0_start_1008_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1008_update_completed_
      -- 
    ack_2071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1008_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block0_start_1011_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_Update/req
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_update_start_
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_sample_completed_
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1011_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block0_start_1011_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	373 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block0_start_1011_update_completed_
      -- 
    ack_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1011_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	234 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_Update/req
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_update_start_
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_Sample/ack
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1014_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block1_start_1014_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_Sample/req
      -- CP-element group 264: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1014_update_completed_
      -- 
    ack_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1014_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block1_start_1017_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_update_start_
      -- CP-element group 265: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_Update/req
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1017_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block1_start_1017_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1017_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_Sample/req
      -- 
    ack_2113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1017_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block1_start_1020_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_update_start_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_Update/req
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1020_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block1_start_1020_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1020_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_Sample/$entry
      -- 
    ack_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1020_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block1_start_1023_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_update_start_
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_Update/req
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_Sample/$exit
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1023_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block1_start_1023_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1023_Update/$exit
      -- 
    ack_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1023_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block1_start_1026_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_Update/req
      -- CP-element group 271: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_update_start_
      -- CP-element group 271: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_sample_completed_
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1026_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block1_start_1026_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1026_update_completed_
      -- 
    ack_2155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1026_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block1_start_1029_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_Update/req
      -- CP-element group 273: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_update_start_
      -- CP-element group 273: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_sample_completed_
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1029_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block1_start_1029_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1029_update_completed_
      -- 
    ack_2169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1029_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block1_start_1032_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_sample_completed_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_Update/req
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_Sample/ack
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1032_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block1_start_1032_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1032_Update/$exit
      -- 
    ack_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1032_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block1_start_1035_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_Update/req
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_update_start_
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_sample_completed_
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1035_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block1_start_1035_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1035_update_completed_
      -- 
    ack_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1035_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block1_start_1038_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_Update/req
      -- CP-element group 279: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_update_start_
      -- CP-element group 279: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_sample_completed_
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1038_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block1_start_1038_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1038_update_completed_
      -- 
    ack_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1038_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	234 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_sample_completed_
      -- 
    ra_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1049_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	234 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1049_update_completed_
      -- 
    ca_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1049_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_sample_start_
      -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block1_start_1051_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(280) & convTranspose_CP_39_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_update_start_
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_Update/req
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1051_inst_ack_0, ack => convTranspose_CP_39_elements(284)); -- 
    req_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_Block1_start_1051_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1051_Update/ack
      -- 
    ack_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1051_inst_ack_1, ack => convTranspose_CP_39_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	234 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_sample_completed_
      -- 
    ra_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1056_inst_ack_0, ack => convTranspose_CP_39_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	234 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1056_update_completed_
      -- 
    ca_2253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1056_inst_ack_1, ack => convTranspose_CP_39_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_sample_start_
      -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block1_start_1058_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(285) & convTranspose_CP_39_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_Update/req
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_sample_completed_
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1058_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block1_start_1058_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1058_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_sample_start_
      -- 
    ack_2267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1058_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_Block1_start_1061_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_Update/req
      -- CP-element group 291: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_update_start_
      -- CP-element group 291: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_sample_completed_
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1061_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_Block1_start_1061_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1061_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_Sample/req
      -- 
    ack_2281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1061_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(292), ack => WPIPE_Block1_start_1064_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_Update/req
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_Sample/ack
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1064_inst_ack_0, ack => convTranspose_CP_39_elements(293)); -- 
    req_2294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block1_start_1064_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1064_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_sample_start_
      -- 
    ack_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1064_inst_ack_1, ack => convTranspose_CP_39_elements(294)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block1_start_1067_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_Update/req
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_sample_completed_
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1067_inst_ack_0, ack => convTranspose_CP_39_elements(295)); -- 
    req_2308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => WPIPE_Block1_start_1067_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	373 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block1_start_1067_update_completed_
      -- 
    ack_2309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1067_inst_ack_1, ack => convTranspose_CP_39_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	234 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_update_start_
      -- CP-element group 297: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_Update/req
      -- CP-element group 297: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_Sample/ack
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1070_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_Block2_start_1070_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1070_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_Sample/$entry
      -- 
    ack_2323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1070_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block2_start_1073_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_update_start_
      -- CP-element group 299: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_Update/req
      -- CP-element group 299: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_Sample/$exit
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1073_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block2_start_1073_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1073_update_completed_
      -- 
    ack_2337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1073_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_Block2_start_1076_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_Update/req
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_sample_completed_
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1076_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    req_2350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block2_start_1076_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1076_Update/ack
      -- 
    ack_2351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1076_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block2_start_1079_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_update_start_
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_Update/req
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1079_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_Block2_start_1079_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1079_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_sample_start_
      -- 
    ack_2365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1079_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block2_start_1082_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_update_start_
      -- CP-element group 305: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_Update/req
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1082_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block2_start_1082_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1082_Update/ack
      -- 
    ack_2379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1082_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(306), ack => WPIPE_Block2_start_1085_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_update_start_
      -- CP-element group 307: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_Update/req
      -- CP-element group 307: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_Update/$entry
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1085_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block2_start_1085_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1085_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_Sample/req
      -- 
    ack_2393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1085_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block2_start_1088_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_update_start_
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_Update/req
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1088_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block2_start_1088_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1088_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_Sample/req
      -- 
    ack_2407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1088_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_Block2_start_1091_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_update_start_
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_Update/req
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1091_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_Block2_start_1091_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1091_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_Sample/req
      -- 
    ack_2421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1091_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(312), ack => WPIPE_Block2_start_1094_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_update_start_
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_Update/req
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1094_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    req_2434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => WPIPE_Block2_start_1094_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1094_Update/ack
      -- 
    ack_2435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1094_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	234 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_Sample/ra
      -- 
    ra_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	234 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1105_Update/ca
      -- 
    ca_2449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	316 
    -- CP-element group 317: 	314 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_Sample/req
      -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_Block2_start_1107_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(316) & convTranspose_CP_39_elements(314);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_update_start_
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_Update/req
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1107_inst_ack_0, ack => convTranspose_CP_39_elements(318)); -- 
    req_2462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(318), ack => WPIPE_Block2_start_1107_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1107_Update/ack
      -- 
    ack_2463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1107_inst_ack_1, ack => convTranspose_CP_39_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	234 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_Sample/ra
      -- 
    ra_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_0, ack => convTranspose_CP_39_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	234 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1112_Update/ca
      -- 
    ca_2477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_1, ack => convTranspose_CP_39_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_Sample/req
      -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => WPIPE_Block2_start_1114_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(319) & convTranspose_CP_39_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_update_start_
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_Update/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1114_inst_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    req_2490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_Block2_start_1114_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1114_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_Sample/req
      -- 
    ack_2491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1114_inst_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_Block2_start_1117_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_update_start_
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_Update/req
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1117_inst_ack_0, ack => convTranspose_CP_39_elements(325)); -- 
    req_2504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => WPIPE_Block2_start_1117_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1117_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_Sample/req
      -- 
    ack_2505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1117_inst_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => WPIPE_Block2_start_1120_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_update_start_
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_Update/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1120_inst_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    req_2518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => WPIPE_Block2_start_1120_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1120_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_Sample/req
      -- 
    ack_2519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1120_inst_ack_1, ack => convTranspose_CP_39_elements(328)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(328), ack => WPIPE_Block2_start_1123_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_update_start_
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_Update/req
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1123_inst_ack_0, ack => convTranspose_CP_39_elements(329)); -- 
    req_2532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(329), ack => WPIPE_Block2_start_1123_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	373 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block2_start_1123_Update/ack
      -- 
    ack_2533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1123_inst_ack_1, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	234 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_update_start_
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_Update/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1126_inst_ack_0, ack => convTranspose_CP_39_elements(331)); -- 
    req_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => WPIPE_Block3_start_1126_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1126_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_Sample/req
      -- 
    ack_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1126_inst_ack_1, ack => convTranspose_CP_39_elements(332)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(332), ack => WPIPE_Block3_start_1129_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_update_start_
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_Update/req
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1129_inst_ack_0, ack => convTranspose_CP_39_elements(333)); -- 
    req_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => WPIPE_Block3_start_1129_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1129_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_Sample/req
      -- 
    ack_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1129_inst_ack_1, ack => convTranspose_CP_39_elements(334)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(334), ack => WPIPE_Block3_start_1132_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_update_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_Update/req
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1132_inst_ack_0, ack => convTranspose_CP_39_elements(335)); -- 
    req_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => WPIPE_Block3_start_1132_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1132_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_Sample/req
      -- 
    ack_2575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1132_inst_ack_1, ack => convTranspose_CP_39_elements(336)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(336), ack => WPIPE_Block3_start_1135_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_update_start_
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_Update/req
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1135_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    req_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => WPIPE_Block3_start_1135_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1135_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_Sample/req
      -- 
    ack_2589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1135_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(338), ack => WPIPE_Block3_start_1138_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_update_start_
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_Update/req
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1138_inst_ack_0, ack => convTranspose_CP_39_elements(339)); -- 
    req_2602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => WPIPE_Block3_start_1138_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1138_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_Sample/req
      -- 
    ack_2603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1138_inst_ack_1, ack => convTranspose_CP_39_elements(340)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(340), ack => WPIPE_Block3_start_1141_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_update_start_
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_Update/req
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1141_inst_ack_0, ack => convTranspose_CP_39_elements(341)); -- 
    req_2616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(341), ack => WPIPE_Block3_start_1141_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1141_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_Sample/req
      -- 
    ack_2617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1141_inst_ack_1, ack => convTranspose_CP_39_elements(342)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(342), ack => WPIPE_Block3_start_1144_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_update_start_
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_Update/req
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1144_inst_ack_0, ack => convTranspose_CP_39_elements(343)); -- 
    req_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_Block3_start_1144_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1144_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_Sample/req
      -- 
    ack_2631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1144_inst_ack_1, ack => convTranspose_CP_39_elements(344)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(344), ack => WPIPE_Block3_start_1147_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_update_start_
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_Update/req
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1147_inst_ack_0, ack => convTranspose_CP_39_elements(345)); -- 
    req_2644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => WPIPE_Block3_start_1147_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1147_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_Sample/req
      -- 
    ack_2645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1147_inst_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => WPIPE_Block3_start_1150_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_update_start_
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_Update/req
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1150_inst_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    req_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(347), ack => WPIPE_Block3_start_1150_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1150_Update/ack
      -- 
    ack_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1150_inst_ack_1, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	234 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_Sample/ra
      -- 
    ra_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1161_inst_ack_0, ack => convTranspose_CP_39_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	234 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1161_Update/ca
      -- 
    ca_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1161_inst_ack_1, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_Sample/req
      -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => WPIPE_Block3_start_1163_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(348) & convTranspose_CP_39_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_update_start_
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_Update/req
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1163_inst_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    req_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_Block3_start_1163_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1163_Update/ack
      -- 
    ack_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1163_inst_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	234 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_Sample/ra
      -- 
    ra_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_0, ack => convTranspose_CP_39_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	234 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/type_cast_1168_Update/ca
      -- 
    ca_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1168_inst_ack_1, ack => convTranspose_CP_39_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_Sample/req
      -- 
    req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(356), ack => WPIPE_Block3_start_1170_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(353) & convTranspose_CP_39_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_update_start_
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_Update/req
      -- 
    ack_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1170_inst_ack_0, ack => convTranspose_CP_39_elements(357)); -- 
    req_2714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(357), ack => WPIPE_Block3_start_1170_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1170_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_Sample/req
      -- 
    ack_2715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1170_inst_ack_1, ack => convTranspose_CP_39_elements(358)); -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(358), ack => WPIPE_Block3_start_1173_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_update_start_
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_Update/req
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1173_inst_ack_0, ack => convTranspose_CP_39_elements(359)); -- 
    req_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => WPIPE_Block3_start_1173_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1173_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_Sample/req
      -- 
    ack_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1173_inst_ack_1, ack => convTranspose_CP_39_elements(360)); -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => WPIPE_Block3_start_1176_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_update_start_
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_Update/req
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1176_inst_ack_0, ack => convTranspose_CP_39_elements(361)); -- 
    req_2742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(361), ack => WPIPE_Block3_start_1176_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1176_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_Sample/req
      -- 
    ack_2743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1176_inst_ack_1, ack => convTranspose_CP_39_elements(362)); -- 
    req_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(362), ack => WPIPE_Block3_start_1179_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_update_start_
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_Update/req
      -- 
    ack_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1179_inst_ack_0, ack => convTranspose_CP_39_elements(363)); -- 
    req_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(363), ack => WPIPE_Block3_start_1179_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	373 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/WPIPE_Block3_start_1179_Update/ack
      -- 
    ack_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1179_inst_ack_1, ack => convTranspose_CP_39_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	234 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_update_start_
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_Sample/ra
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_Update/cr
      -- 
    ra_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1183_inst_ack_0, ack => convTranspose_CP_39_elements(365)); -- 
    cr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(365), ack => RPIPE_Block0_done_1183_inst_req_1); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	373 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block0_done_1183_Update/ca
      -- 
    ca_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1183_inst_ack_1, ack => convTranspose_CP_39_elements(366)); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	234 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_update_start_
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_Sample/ra
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_Update/cr
      -- 
    ra_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1186_inst_ack_0, ack => convTranspose_CP_39_elements(367)); -- 
    cr_2784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => RPIPE_Block1_done_1186_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	373 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block1_done_1186_Update/ca
      -- 
    ca_2785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1186_inst_ack_1, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	234 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_update_start_
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_Sample/ra
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_Update/cr
      -- 
    ra_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1189_inst_ack_0, ack => convTranspose_CP_39_elements(369)); -- 
    cr_2798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(369), ack => RPIPE_Block2_done_1189_inst_req_1); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	373 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block2_done_1189_Update/ca
      -- 
    ca_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1189_inst_ack_1, ack => convTranspose_CP_39_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	234 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_update_start_
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_Sample/ra
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_Update/cr
      -- 
    ra_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1192_inst_ack_0, ack => convTranspose_CP_39_elements(371)); -- 
    cr_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => RPIPE_Block3_done_1192_inst_req_1); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/RPIPE_Block3_done_1192_Update/ca
      -- 
    ca_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1192_inst_ack_1, ack => convTranspose_CP_39_elements(372)); -- 
    -- CP-element group 373:  join  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	330 
    -- CP-element group 373: 	364 
    -- CP-element group 373: 	366 
    -- CP-element group 373: 	368 
    -- CP-element group 373: 	370 
    -- CP-element group 373: 	372 
    -- CP-element group 373: 	262 
    -- CP-element group 373: 	296 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	377 
    -- CP-element group 373: 	379 
    -- CP-element group 373: 	381 
    -- CP-element group 373: 	383 
    -- CP-element group 373: 	385 
    -- CP-element group 373: 	387 
    -- CP-element group 373: 	389 
    -- CP-element group 373: 	391 
    -- CP-element group 373: 	393 
    -- CP-element group 373:  members (37) 
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193__exit__
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304__entry__
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_972_to_assign_stmt_1193/$exit
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_Sample/crr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_Update/ccr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_Update/cr
      -- 
    crr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1196_call_req_0); -- 
    ccr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1196_call_req_1); -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1200_inst_req_1); -- 
    cr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1209_inst_req_1); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1219_inst_req_1); -- 
    cr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1229_inst_req_1); -- 
    cr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1239_inst_req_1); -- 
    cr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1249_inst_req_1); -- 
    cr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1259_inst_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1269_inst_req_1); -- 
    cr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1279_inst_req_1); -- 
    convTranspose_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(330) & convTranspose_CP_39_elements(364) & convTranspose_CP_39_elements(366) & convTranspose_CP_39_elements(368) & convTranspose_CP_39_elements(370) & convTranspose_CP_39_elements(372) & convTranspose_CP_39_elements(262) & convTranspose_CP_39_elements(296);
      gj_convTranspose_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_Sample/cra
      -- 
    cra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1196_call_ack_0, ack => convTranspose_CP_39_elements(374)); -- 
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/call_stmt_1196_Update/cca
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_Sample/rr
      -- 
    cca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1196_call_ack_1, ack => convTranspose_CP_39_elements(375)); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => type_cast_1200_inst_req_0); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_Sample/ra
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1200_inst_ack_0, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  fork  transition  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	373 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377: 	380 
    -- CP-element group 377: 	382 
    -- CP-element group 377: 	384 
    -- CP-element group 377: 	386 
    -- CP-element group 377: 	388 
    -- CP-element group 377: 	390 
    -- CP-element group 377: 	392 
    -- CP-element group 377:  members (27) 
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1200_Update/ca
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_Sample/rr
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1200_inst_ack_1, ack => convTranspose_CP_39_elements(377)); -- 
    rr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1209_inst_req_0); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1219_inst_req_0); -- 
    rr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1229_inst_req_0); -- 
    rr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1239_inst_req_0); -- 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1249_inst_req_0); -- 
    rr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1259_inst_req_0); -- 
    rr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1269_inst_req_0); -- 
    rr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1279_inst_req_0); -- 
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_Sample/ra
      -- 
    ra_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1209_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	373 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	414 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1209_Update/ca
      -- 
    ca_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1209_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	377 
    -- CP-element group 380: successors 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_Sample/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1219_inst_ack_0, ack => convTranspose_CP_39_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	373 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	411 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1219_Update/ca
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1219_inst_ack_1, ack => convTranspose_CP_39_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	377 
    -- CP-element group 382: successors 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_Sample/ra
      -- 
    ra_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1229_inst_ack_0, ack => convTranspose_CP_39_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	373 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	408 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1229_Update/ca
      -- 
    ca_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1229_inst_ack_1, ack => convTranspose_CP_39_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	377 
    -- CP-element group 384: successors 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_Sample/ra
      -- 
    ra_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	373 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	405 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1239_Update/ca
      -- 
    ca_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	377 
    -- CP-element group 386: successors 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_Sample/ra
      -- 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1249_inst_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	373 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	402 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1249_Update/ca
      -- 
    ca_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1249_inst_ack_1, ack => convTranspose_CP_39_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	377 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_sample_completed_
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_Sample/ra
      -- 
    ra_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_0, ack => convTranspose_CP_39_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	373 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	399 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1259_Update/ca
      -- 
    ca_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_1, ack => convTranspose_CP_39_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	377 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_Sample/ra
      -- 
    ra_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	373 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	396 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1269_Update/ca
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1269_inst_ack_1, ack => convTranspose_CP_39_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	377 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_Sample/ra
      -- 
    ra_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_0, ack => convTranspose_CP_39_elements(392)); -- 
    -- CP-element group 393:  transition  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	373 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (6) 
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/type_cast_1279_Update/ca
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_Sample/req
      -- 
    ca_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_1, ack => convTranspose_CP_39_elements(393)); -- 
    req_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(393), ack => WPIPE_ConvTranspose_output_pipe_1281_inst_req_0); -- 
    -- CP-element group 394:  transition  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (6) 
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_Update/req
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_update_start_
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_Sample/ack
      -- 
    ack_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0, ack => convTranspose_CP_39_elements(394)); -- 
    req_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(394), ack => WPIPE_ConvTranspose_output_pipe_1281_inst_req_1); -- 
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_Update/ack
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1281_update_completed_
      -- 
    ack_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1, ack => convTranspose_CP_39_elements(395)); -- 
    -- CP-element group 396:  join  transition  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	391 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_Sample/req
      -- 
    req_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(396), ack => WPIPE_ConvTranspose_output_pipe_1284_inst_req_0); -- 
    convTranspose_cp_element_group_396: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_396"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(391) & convTranspose_CP_39_elements(395);
      gj_convTranspose_cp_element_group_396 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(396), clk => clk, reset => reset); --
    end block;
    -- CP-element group 397:  transition  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (6) 
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_update_start_
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_Update/req
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_sample_completed_
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_Sample/ack
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_Sample/$exit
      -- 
    ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0, ack => convTranspose_CP_39_elements(397)); -- 
    req_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => WPIPE_ConvTranspose_output_pipe_1284_inst_req_1); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_Update/$exit
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_Update/ack
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1284_update_completed_
      -- 
    ack_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1, ack => convTranspose_CP_39_elements(398)); -- 
    -- CP-element group 399:  join  transition  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	389 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_sample_start_
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_Sample/$entry
      -- 
    req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(399), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_0); -- 
    convTranspose_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(389) & convTranspose_CP_39_elements(398);
      gj_convTranspose_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  transition  input  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (6) 
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_sample_completed_
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_update_start_
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_Update/req
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_Sample/ack
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_Sample/$exit
      -- 
    ack_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0, ack => convTranspose_CP_39_elements(400)); -- 
    req_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(400), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_1); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_update_completed_
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_Update/ack
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1287_Update/$exit
      -- 
    ack_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1, ack => convTranspose_CP_39_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	387 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_Sample/req
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_Sample/$entry
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_sample_start_
      -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_0); -- 
    convTranspose_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(387) & convTranspose_CP_39_elements(401);
      gj_convTranspose_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  transition  input  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (6) 
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_Update/req
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_Sample/ack
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_update_start_
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_sample_completed_
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0, ack => convTranspose_CP_39_elements(403)); -- 
    req_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(403), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_1); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_Update/ack
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1290_update_completed_
      -- 
    ack_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1, ack => convTranspose_CP_39_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	385 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_Sample/req
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_sample_start_
      -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(405), ack => WPIPE_ConvTranspose_output_pipe_1293_inst_req_0); -- 
    convTranspose_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(385) & convTranspose_CP_39_elements(404);
      gj_convTranspose_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (6) 
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_Update/req
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_Sample/ack
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_Sample/$exit
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_update_start_
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_sample_completed_
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0, ack => convTranspose_CP_39_elements(406)); -- 
    req_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => WPIPE_ConvTranspose_output_pipe_1293_inst_req_1); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_Update/ack
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_Update/$exit
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1293_update_completed_
      -- 
    ack_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1, ack => convTranspose_CP_39_elements(407)); -- 
    -- CP-element group 408:  join  transition  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	383 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_Sample/req
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_sample_start_
      -- 
    req_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(408), ack => WPIPE_ConvTranspose_output_pipe_1296_inst_req_0); -- 
    convTranspose_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(383) & convTranspose_CP_39_elements(407);
      gj_convTranspose_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  transition  input  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (6) 
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_Update/req
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_Update/$entry
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_Sample/ack
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_update_start_
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_sample_completed_
      -- 
    ack_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0, ack => convTranspose_CP_39_elements(409)); -- 
    req_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(409), ack => WPIPE_ConvTranspose_output_pipe_1296_inst_req_1); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_Update/ack
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1296_update_completed_
      -- 
    ack_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1, ack => convTranspose_CP_39_elements(410)); -- 
    -- CP-element group 411:  join  transition  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	381 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_Sample/req
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_sample_start_
      -- 
    req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => WPIPE_ConvTranspose_output_pipe_1299_inst_req_0); -- 
    convTranspose_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(381) & convTranspose_CP_39_elements(410);
      gj_convTranspose_cp_element_group_411 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_update_start_
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_Update/req
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_Sample/ack
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_sample_completed_
      -- 
    ack_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0, ack => convTranspose_CP_39_elements(412)); -- 
    req_3053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(412), ack => WPIPE_ConvTranspose_output_pipe_1299_inst_req_1); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_Update/ack
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_update_completed_
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1299_Update/$exit
      -- 
    ack_3054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1, ack => convTranspose_CP_39_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	379 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_sample_start_
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_Sample/req
      -- 
    req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(414), ack => WPIPE_ConvTranspose_output_pipe_1302_inst_req_0); -- 
    convTranspose_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(379) & convTranspose_CP_39_elements(413);
      gj_convTranspose_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_update_start_
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_sample_completed_
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_Update/req
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_Update/$entry
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_Sample/ack
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_Sample/$exit
      -- 
    ack_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0, ack => convTranspose_CP_39_elements(415)); -- 
    req_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(415), ack => WPIPE_ConvTranspose_output_pipe_1302_inst_req_1); -- 
    -- CP-element group 416:  branch  transition  place  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416: 	418 
    -- CP-element group 416:  members (13) 
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304__exit__
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1306__entry__
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_update_completed_
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1306_else_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1306_if_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1306_eval_test/branch_req
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1306_eval_test/$exit
      -- CP-element group 416: 	 branch_block_stmt_32/R_cmp264505_1307_place
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1306_eval_test/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1306_dead_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_Update/ack
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/WPIPE_ConvTranspose_output_pipe_1302_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1196_to_assign_stmt_1304/$exit
      -- 
    ack_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1, ack => convTranspose_CP_39_elements(416)); -- 
    branch_req_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(416), ack => if_stmt_1306_branch_req_0); -- 
    -- CP-element group 417:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	419 
    -- CP-element group 417: 	420 
    -- CP-element group 417:  members (18) 
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1312__exit__
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347__entry__
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_Update/cr
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_Sample/rr
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_update_start_
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_sample_start_
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/forx_xend273_bbx_xnph
      -- CP-element group 417: 	 branch_block_stmt_32/if_stmt_1306_if_link/if_choice_transition
      -- CP-element group 417: 	 branch_block_stmt_32/if_stmt_1306_if_link/$exit
      -- CP-element group 417: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1312_PhiReqMerge
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1312_PhiAck/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1312_PhiAck/$exit
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1312_PhiAck/dummy
      -- 
    if_choice_transition_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1306_branch_ack_1, ack => convTranspose_CP_39_elements(417)); -- 
    cr_3103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => type_cast_1333_inst_req_1); -- 
    rr_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => type_cast_1333_inst_req_0); -- 
    -- CP-element group 418:  transition  place  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	416 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	496 
    -- CP-element group 418:  members (5) 
      -- CP-element group 418: 	 branch_block_stmt_32/forx_xend273_forx_xend500
      -- CP-element group 418: 	 branch_block_stmt_32/if_stmt_1306_else_link/else_choice_transition
      -- CP-element group 418: 	 branch_block_stmt_32/if_stmt_1306_else_link/$exit
      -- CP-element group 418: 	 branch_block_stmt_32/forx_xend273_forx_xend500_PhiReq/$entry
      -- CP-element group 418: 	 branch_block_stmt_32/forx_xend273_forx_xend500_PhiReq/$exit
      -- 
    else_choice_transition_3085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1306_branch_ack_0, ack => convTranspose_CP_39_elements(418)); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: successors 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_Sample/ra
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_sample_completed_
      -- 
    ra_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1333_inst_ack_0, ack => convTranspose_CP_39_elements(419)); -- 
    -- CP-element group 420:  transition  place  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	417 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	490 
    -- CP-element group 420:  members (9) 
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347__exit__
      -- CP-element group 420: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_Update/ca
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/type_cast_1333_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1318_to_assign_stmt_1347/$exit
      -- CP-element group 420: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/$entry
      -- CP-element group 420: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1350/$entry
      -- CP-element group 420: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/$entry
      -- 
    ca_3104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1333_inst_ack_1, ack => convTranspose_CP_39_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	495 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	466 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_sample_complete
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_Sample/ack
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_Sample/$exit
      -- 
    ack_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1362_index_offset_ack_0, ack => convTranspose_CP_39_elements(421)); -- 
    -- CP-element group 422:  transition  input  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	495 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (11) 
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_Update/$exit
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_Update/ack
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_base_plus_offset/$entry
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_offset_calculated
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_root_address_calculated
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_sample_start_
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_request/req
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_request/$entry
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_base_plus_offset/sum_rename_ack
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_base_plus_offset/sum_rename_req
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_base_plus_offset/$exit
      -- 
    ack_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1362_index_offset_ack_1, ack => convTranspose_CP_39_elements(422)); -- 
    req_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(422), ack => addr_of_1363_final_reg_req_0); -- 
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_sample_completed_
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_request/ack
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_request/$exit
      -- 
    ack_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1363_final_reg_ack_0, ack => convTranspose_CP_39_elements(423)); -- 
    -- CP-element group 424:  join  fork  transition  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	495 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (24) 
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_update_completed_
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_word_addrgen/root_register_ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_word_addrgen/root_register_req
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_word_addrgen/$exit
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_word_addrgen/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_plus_offset/sum_rename_ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_plus_offset/sum_rename_req
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_plus_offset/$exit
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_plus_offset/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_addr_resize/base_resize_ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_addr_resize/base_resize_req
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_addr_resize/$exit
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_addr_resize/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_address_resized
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_base_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_complete/ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_complete/$exit
      -- 
    ack_3153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1363_final_reg_ack_1, ack => convTranspose_CP_39_elements(424)); -- 
    rr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => ptr_deref_1367_load_0_req_0); -- 
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425:  members (5) 
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Sample/word_access_start/word_0/ra
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Sample/word_access_start/word_0/$exit
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Sample/word_access_start/$exit
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_sample_completed_
      -- 
    ra_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1367_load_0_ack_0, ack => convTranspose_CP_39_elements(425)); -- 
    -- CP-element group 426:  fork  transition  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	495 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426: 	429 
    -- CP-element group 426: 	431 
    -- CP-element group 426: 	433 
    -- CP-element group 426: 	435 
    -- CP-element group 426: 	437 
    -- CP-element group 426: 	439 
    -- CP-element group 426: 	441 
    -- CP-element group 426:  members (33) 
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/ptr_deref_1367_Merge/merge_ack
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/ptr_deref_1367_Merge/merge_req
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/ptr_deref_1367_Merge/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/ptr_deref_1367_Merge/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/word_access_complete/word_0/ca
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/word_access_complete/word_0/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/word_access_complete/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_update_completed_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_Sample/$entry
      -- 
    ca_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1367_load_0_ack_1, ack => convTranspose_CP_39_elements(426)); -- 
    rr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1371_inst_req_0); -- 
    rr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1381_inst_req_0); -- 
    rr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1391_inst_req_0); -- 
    rr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1401_inst_req_0); -- 
    rr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1411_inst_req_0); -- 
    rr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1421_inst_req_0); -- 
    rr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1431_inst_req_0); -- 
    rr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1441_inst_req_0); -- 
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_Sample/$exit
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_Sample/ra
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_sample_completed_
      -- 
    ra_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_0, ack => convTranspose_CP_39_elements(427)); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	495 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	463 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_Update/ca
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_update_completed_
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_Update/$exit
      -- 
    ca_3217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_1, ack => convTranspose_CP_39_elements(428)); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	426 
    -- CP-element group 429: successors 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_sample_completed_
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_Sample/$exit
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_Sample/ra
      -- 
    ra_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1381_inst_ack_0, ack => convTranspose_CP_39_elements(429)); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	495 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	460 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_update_completed_
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_Update/ca
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_Update/$exit
      -- 
    ca_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1381_inst_ack_1, ack => convTranspose_CP_39_elements(430)); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	426 
    -- CP-element group 431: successors 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_Sample/ra
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_sample_completed_
      -- 
    ra_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_0, ack => convTranspose_CP_39_elements(431)); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	495 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	457 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_Update/ca
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_update_completed_
      -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_1, ack => convTranspose_CP_39_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	426 
    -- CP-element group 433: successors 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_Sample/ra
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_Sample/$exit
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_sample_completed_
      -- 
    ra_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1401_inst_ack_0, ack => convTranspose_CP_39_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	495 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	454 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_Update/ca
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_Update/$exit
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_update_completed_
      -- 
    ca_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1401_inst_ack_1, ack => convTranspose_CP_39_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	426 
    -- CP-element group 435: successors 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_sample_completed_
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_Sample/ra
      -- 
    ra_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_0, ack => convTranspose_CP_39_elements(435)); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	495 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	451 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_update_completed_
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_Update/ca
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_Update/$exit
      -- 
    ca_3273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_1, ack => convTranspose_CP_39_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	426 
    -- CP-element group 437: successors 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_Sample/ra
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_Sample/$exit
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_sample_completed_
      -- 
    ra_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1421_inst_ack_0, ack => convTranspose_CP_39_elements(437)); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	495 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	448 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_Update/ca
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_Update/$exit
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_update_completed_
      -- 
    ca_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1421_inst_ack_1, ack => convTranspose_CP_39_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	426 
    -- CP-element group 439: successors 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_Sample/ra
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_Sample/$exit
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_sample_completed_
      -- 
    ra_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1431_inst_ack_0, ack => convTranspose_CP_39_elements(439)); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	495 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	445 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_Update/$exit
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_Update/ca
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_update_completed_
      -- 
    ca_3301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1431_inst_ack_1, ack => convTranspose_CP_39_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	426 
    -- CP-element group 441: successors 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_sample_completed_
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_Sample/ra
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_Sample/$exit
      -- 
    ra_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1441_inst_ack_0, ack => convTranspose_CP_39_elements(441)); -- 
    -- CP-element group 442:  transition  input  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	495 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442:  members (6) 
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_Update/ca
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_Update/$exit
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_Sample/req
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_Sample/$entry
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_sample_start_
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_update_completed_
      -- 
    ca_3315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1441_inst_ack_1, ack => convTranspose_CP_39_elements(442)); -- 
    req_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(442), ack => WPIPE_ConvTranspose_output_pipe_1443_inst_req_0); -- 
    -- CP-element group 443:  transition  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (6) 
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_Update/req
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_Sample/ack
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_update_start_
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_sample_completed_
      -- 
    ack_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1443_inst_ack_0, ack => convTranspose_CP_39_elements(443)); -- 
    req_3328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(443), ack => WPIPE_ConvTranspose_output_pipe_1443_inst_req_1); -- 
    -- CP-element group 444:  transition  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_Update/ack
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1443_update_completed_
      -- 
    ack_3329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1443_inst_ack_1, ack => convTranspose_CP_39_elements(444)); -- 
    -- CP-element group 445:  join  transition  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	440 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_Sample/req
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_sample_start_
      -- 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => WPIPE_ConvTranspose_output_pipe_1446_inst_req_0); -- 
    convTranspose_cp_element_group_445: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_445"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(440) & convTranspose_CP_39_elements(444);
      gj_convTranspose_cp_element_group_445 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(445), clk => clk, reset => reset); --
    end block;
    -- CP-element group 446:  transition  input  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (6) 
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_Update/req
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_Sample/ack
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_Sample/$exit
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_update_start_
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_sample_completed_
      -- 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1446_inst_ack_0, ack => convTranspose_CP_39_elements(446)); -- 
    req_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(446), ack => WPIPE_ConvTranspose_output_pipe_1446_inst_req_1); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_Update/ack
      -- CP-element group 447: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_Update/$exit
      -- CP-element group 447: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1446_update_completed_
      -- 
    ack_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1446_inst_ack_1, ack => convTranspose_CP_39_elements(447)); -- 
    -- CP-element group 448:  join  transition  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	438 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_Sample/$entry
      -- CP-element group 448: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_sample_start_
      -- CP-element group 448: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_Sample/req
      -- 
    req_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(448), ack => WPIPE_ConvTranspose_output_pipe_1449_inst_req_0); -- 
    convTranspose_cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(438) & convTranspose_CP_39_elements(447);
      gj_convTranspose_cp_element_group_448 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 449:  transition  input  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (6) 
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_sample_completed_
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_Update/req
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_update_start_
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_Sample/ack
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_Sample/$exit
      -- 
    ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0, ack => convTranspose_CP_39_elements(449)); -- 
    req_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(449), ack => WPIPE_ConvTranspose_output_pipe_1449_inst_req_1); -- 
    -- CP-element group 450:  transition  input  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_Update/ack
      -- CP-element group 450: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_update_completed_
      -- CP-element group 450: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1449_Update/$exit
      -- 
    ack_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1, ack => convTranspose_CP_39_elements(450)); -- 
    -- CP-element group 451:  join  transition  output  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	436 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_Sample/req
      -- CP-element group 451: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_sample_start_
      -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(451), ack => WPIPE_ConvTranspose_output_pipe_1452_inst_req_0); -- 
    convTranspose_cp_element_group_451: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_451"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(436) & convTranspose_CP_39_elements(450);
      gj_convTranspose_cp_element_group_451 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(451), clk => clk, reset => reset); --
    end block;
    -- CP-element group 452:  transition  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (6) 
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_Update/req
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_Sample/ack
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_update_start_
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_sample_completed_
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0, ack => convTranspose_CP_39_elements(452)); -- 
    req_3370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => WPIPE_ConvTranspose_output_pipe_1452_inst_req_1); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_Update/ack
      -- CP-element group 453: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1452_update_completed_
      -- 
    ack_3371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1, ack => convTranspose_CP_39_elements(453)); -- 
    -- CP-element group 454:  join  transition  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	434 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_sample_start_
      -- CP-element group 454: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_Sample/req
      -- 
    req_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(454), ack => WPIPE_ConvTranspose_output_pipe_1455_inst_req_0); -- 
    convTranspose_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(434) & convTranspose_CP_39_elements(453);
      gj_convTranspose_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  transition  input  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (6) 
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_sample_completed_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_Sample/ack
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_Update/req
      -- 
    ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0, ack => convTranspose_CP_39_elements(455)); -- 
    req_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => WPIPE_ConvTranspose_output_pipe_1455_inst_req_1); -- 
    -- CP-element group 456:  transition  input  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_update_completed_
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1455_Update/ack
      -- 
    ack_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1, ack => convTranspose_CP_39_elements(456)); -- 
    -- CP-element group 457:  join  transition  output  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	432 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_sample_start_
      -- CP-element group 457: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_Sample/$entry
      -- CP-element group 457: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_Sample/req
      -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(457), ack => WPIPE_ConvTranspose_output_pipe_1458_inst_req_0); -- 
    convTranspose_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(432) & convTranspose_CP_39_elements(456);
      gj_convTranspose_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  transition  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (6) 
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_sample_completed_
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_update_start_
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_Sample/$exit
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_Sample/ack
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_Update/req
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0, ack => convTranspose_CP_39_elements(458)); -- 
    req_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => WPIPE_ConvTranspose_output_pipe_1458_inst_req_1); -- 
    -- CP-element group 459:  transition  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_update_completed_
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_Update/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1458_Update/ack
      -- 
    ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1, ack => convTranspose_CP_39_elements(459)); -- 
    -- CP-element group 460:  join  transition  output  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	430 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_sample_start_
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_Sample/req
      -- 
    req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(460), ack => WPIPE_ConvTranspose_output_pipe_1461_inst_req_0); -- 
    convTranspose_cp_element_group_460: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_460"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(430) & convTranspose_CP_39_elements(459);
      gj_convTranspose_cp_element_group_460 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(460), clk => clk, reset => reset); --
    end block;
    -- CP-element group 461:  transition  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (6) 
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_sample_completed_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_Sample/$exit
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_Sample/ack
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_Update/req
      -- 
    ack_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0, ack => convTranspose_CP_39_elements(461)); -- 
    req_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => WPIPE_ConvTranspose_output_pipe_1461_inst_req_1); -- 
    -- CP-element group 462:  transition  input  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_update_completed_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1461_Update/ack
      -- 
    ack_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1, ack => convTranspose_CP_39_elements(462)); -- 
    -- CP-element group 463:  join  transition  output  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	428 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_Sample/$entry
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_Sample/req
      -- 
    req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(463), ack => WPIPE_ConvTranspose_output_pipe_1464_inst_req_0); -- 
    convTranspose_cp_element_group_463: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_463"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(428) & convTranspose_CP_39_elements(462);
      gj_convTranspose_cp_element_group_463 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(463), clk => clk, reset => reset); --
    end block;
    -- CP-element group 464:  transition  input  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464:  members (6) 
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_update_start_
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_Sample/ack
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_Update/$entry
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_Update/req
      -- 
    ack_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0, ack => convTranspose_CP_39_elements(464)); -- 
    req_3426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(464), ack => WPIPE_ConvTranspose_output_pipe_1464_inst_req_1); -- 
    -- CP-element group 465:  transition  input  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/WPIPE_ConvTranspose_output_pipe_1464_Update/ack
      -- 
    ack_3427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1, ack => convTranspose_CP_39_elements(465)); -- 
    -- CP-element group 466:  branch  join  transition  place  output  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	421 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466: 	468 
    -- CP-element group 466:  members (10) 
      -- CP-element group 466: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477__exit__
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1478__entry__
      -- CP-element group 466: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1478_dead_link/$entry
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1478_eval_test/$entry
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1478_eval_test/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1478_eval_test/branch_req
      -- CP-element group 466: 	 branch_block_stmt_32/R_exitcond1_1479_place
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1478_if_link/$entry
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1478_else_link/$entry
      -- 
    branch_req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(466), ack => if_stmt_1478_branch_req_0); -- 
    convTranspose_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(421) & convTranspose_CP_39_elements(465);
      gj_convTranspose_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  merge  transition  place  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	496 
    -- CP-element group 467:  members (13) 
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1484__exit__
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xend500x_xloopexit_forx_xend500
      -- CP-element group 467: 	 branch_block_stmt_32/if_stmt_1478_if_link/$exit
      -- CP-element group 467: 	 branch_block_stmt_32/if_stmt_1478_if_link/if_choice_transition
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xbody427_forx_xend500x_xloopexit
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$entry
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$exit
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1484_PhiReqMerge
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1484_PhiAck/$entry
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1484_PhiAck/$exit
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1484_PhiAck/dummy
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xend500x_xloopexit_forx_xend500_PhiReq/$entry
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xend500x_xloopexit_forx_xend500_PhiReq/$exit
      -- 
    if_choice_transition_3440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1478_branch_ack_1, ack => convTranspose_CP_39_elements(467)); -- 
    -- CP-element group 468:  fork  transition  place  input  output  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	466 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	491 
    -- CP-element group 468: 	492 
    -- CP-element group 468:  members (12) 
      -- CP-element group 468: 	 branch_block_stmt_32/if_stmt_1478_else_link/$exit
      -- CP-element group 468: 	 branch_block_stmt_32/if_stmt_1478_else_link/else_choice_transition
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/Sample/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/Sample/rr
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/Update/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1478_branch_ack_0, ack => convTranspose_CP_39_elements(468)); -- 
    rr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => type_cast_1356_inst_req_0); -- 
    cr_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => type_cast_1356_inst_req_1); -- 
    -- CP-element group 469:  merge  branch  transition  place  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	165 
    -- CP-element group 469: 	120 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	121 
    -- CP-element group 469: 	122 
    -- CP-element group 469:  members (17) 
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424__exit__
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_430__entry__
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_430__exit__
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431__entry__
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_430/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_430/$exit
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_dead_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_eval_test/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_eval_test/$exit
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_eval_test/branch_req
      -- CP-element group 469: 	 branch_block_stmt_32/R_cmp194509_432_place
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_if_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_else_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424_PhiReqMerge
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/$exit
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/dummy
      -- 
    branch_req_927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => if_stmt_431_branch_req_0); -- 
    convTranspose_CP_39_elements(469) <= OrReduce(convTranspose_CP_39_elements(165) & convTranspose_CP_39_elements(120));
    -- CP-element group 470:  transition  output  delay-element  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	124 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	474 
    -- CP-element group 470:  members (5) 
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_473_konst_delay_trans
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_req
      -- 
    phi_stmt_469_req_3492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_469_req_3492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(470), ack => phi_stmt_469_req_0); -- 
    -- Element group convTranspose_CP_39_elements(470) is a control-delay.
    cp_element_470_delay: control_delay_element  generic map(name => " 470_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(124), ack => convTranspose_CP_39_elements(470), clk => clk, reset =>reset);
    -- CP-element group 471:  transition  input  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	166 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	473 
    -- CP-element group 471:  members (2) 
      -- CP-element group 471: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/$exit
      -- CP-element group 471: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/ra
      -- 
    ra_3512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_475_inst_ack_0, ack => convTranspose_CP_39_elements(471)); -- 
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	166 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472:  members (2) 
      -- CP-element group 472: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/$exit
      -- CP-element group 472: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/ca
      -- 
    ca_3517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_475_inst_ack_1, ack => convTranspose_CP_39_elements(472)); -- 
    -- CP-element group 473:  join  transition  output  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	471 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (6) 
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_req
      -- 
    phi_stmt_469_req_3518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_469_req_3518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(473), ack => phi_stmt_469_req_1); -- 
    convTranspose_cp_element_group_473: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_473"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(471) & convTranspose_CP_39_elements(472);
      gj_convTranspose_cp_element_group_473 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(473), clk => clk, reset => reset); --
    end block;
    -- CP-element group 474:  merge  transition  place  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	470 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (2) 
      -- CP-element group 474: 	 branch_block_stmt_32/merge_stmt_468_PhiReqMerge
      -- CP-element group 474: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(474) <= OrReduce(convTranspose_CP_39_elements(470) & convTranspose_CP_39_elements(473));
    -- CP-element group 475:  fork  transition  place  input  output  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	160 
    -- CP-element group 475: 	163 
    -- CP-element group 475: 	125 
    -- CP-element group 475: 	126 
    -- CP-element group 475: 	128 
    -- CP-element group 475: 	129 
    -- CP-element group 475: 	132 
    -- CP-element group 475: 	136 
    -- CP-element group 475: 	140 
    -- CP-element group 475: 	144 
    -- CP-element group 475: 	148 
    -- CP-element group 475: 	152 
    -- CP-element group 475: 	156 
    -- CP-element group 475:  members (56) 
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_468__exit__
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631__entry__
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resized_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scaled_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_computed_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/index_resize_req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/index_resize_ack
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/scale_rename_req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/scale_rename_ack
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_update_start
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/rr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/phi_stmt_469_ack
      -- 
    phi_stmt_469_ack_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_469_ack_0, ack => convTranspose_CP_39_elements(475)); -- 
    cr_1115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_538_inst_req_1); -- 
    cr_1171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_574_inst_req_1); -- 
    cr_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => ptr_deref_618_store_0_req_1); -- 
    cr_1227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_610_inst_req_1); -- 
    cr_1143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_556_inst_req_1); -- 
    cr_1199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_592_inst_req_1); -- 
    req_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => array_obj_ref_481_index_offset_req_0); -- 
    req_988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => array_obj_ref_481_index_offset_req_1); -- 
    req_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => addr_of_482_final_reg_req_1); -- 
    rr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => RPIPE_ConvTranspose_input_pipe_485_inst_req_0); -- 
    cr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_489_inst_req_1); -- 
    cr_1059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_502_inst_req_1); -- 
    cr_1087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_520_inst_req_1); -- 
    -- CP-element group 476:  transition  output  delay-element  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	168 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	480 
    -- CP-element group 476:  members (5) 
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_682_konst_delay_trans
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_req
      -- 
    phi_stmt_676_req_3546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_req_3546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(476), ack => phi_stmt_676_req_1); -- 
    -- Element group convTranspose_CP_39_elements(476) is a control-delay.
    cp_element_476_delay: control_delay_element  generic map(name => " 476_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(168), ack => convTranspose_CP_39_elements(476), clk => clk, reset =>reset);
    -- CP-element group 477:  transition  input  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	210 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	479 
    -- CP-element group 477:  members (2) 
      -- CP-element group 477: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/$exit
      -- CP-element group 477: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/ra
      -- 
    ra_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_0, ack => convTranspose_CP_39_elements(477)); -- 
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	210 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	479 
    -- CP-element group 478:  members (2) 
      -- CP-element group 478: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/$exit
      -- CP-element group 478: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/ca
      -- 
    ca_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_1, ack => convTranspose_CP_39_elements(478)); -- 
    -- CP-element group 479:  join  transition  output  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	477 
    -- CP-element group 479: 	478 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (6) 
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_req
      -- 
    phi_stmt_676_req_3572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_req_3572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(479), ack => phi_stmt_676_req_0); -- 
    convTranspose_cp_element_group_479: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_479"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(477) & convTranspose_CP_39_elements(478);
      gj_convTranspose_cp_element_group_479 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(479), clk => clk, reset => reset); --
    end block;
    -- CP-element group 480:  merge  transition  place  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	476 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480:  members (2) 
      -- CP-element group 480: 	 branch_block_stmt_32/merge_stmt_675_PhiReqMerge
      -- CP-element group 480: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(480) <= OrReduce(convTranspose_CP_39_elements(476) & convTranspose_CP_39_elements(479));
    -- CP-element group 481:  fork  transition  place  input  output  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	180 
    -- CP-element group 481: 	184 
    -- CP-element group 481: 	188 
    -- CP-element group 481: 	192 
    -- CP-element group 481: 	196 
    -- CP-element group 481: 	176 
    -- CP-element group 481: 	200 
    -- CP-element group 481: 	204 
    -- CP-element group 481: 	207 
    -- CP-element group 481: 	169 
    -- CP-element group 481: 	170 
    -- CP-element group 481: 	172 
    -- CP-element group 481: 	173 
    -- CP-element group 481:  members (56) 
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/merge_stmt_675__exit__
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838__entry__
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/rr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_sample_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scaled_1
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resized_1
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_update_start
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/scale_rename_ack
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/scale_rename_req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/$exit
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/index_resize_ack
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/index_resize_req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/$exit
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_computed_1
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/cr
      -- CP-element group 481: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/$exit
      -- CP-element group 481: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/phi_stmt_676_ack
      -- 
    phi_stmt_676_ack_3577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_676_ack_0, ack => convTranspose_CP_39_elements(481)); -- 
    rr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => RPIPE_ConvTranspose_input_pipe_692_inst_req_0); -- 
    req_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => addr_of_689_final_reg_req_1); -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_727_inst_req_1); -- 
    req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => array_obj_ref_688_index_offset_req_1); -- 
    cr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_696_inst_req_1); -- 
    req_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => array_obj_ref_688_index_offset_req_0); -- 
    cr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_709_inst_req_1); -- 
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_745_inst_req_1); -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_763_inst_req_1); -- 
    cr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_781_inst_req_1); -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_799_inst_req_1); -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_817_inst_req_1); -- 
    cr_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => ptr_deref_825_store_0_req_1); -- 
    -- CP-element group 482:  merge  fork  transition  place  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	209 
    -- CP-element group 482: 	122 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	211 
    -- CP-element group 482: 	212 
    -- CP-element group 482: 	213 
    -- CP-element group 482: 	214 
    -- CP-element group 482: 	215 
    -- CP-element group 482: 	216 
    -- CP-element group 482:  members (25) 
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847__exit__
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875__entry__
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_update_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_update_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_update_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847_PhiReqMerge
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/$exit
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/dummy
      -- 
    rr_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_850_inst_req_0); -- 
    cr_1672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_850_inst_req_1); -- 
    rr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_854_inst_req_0); -- 
    cr_1686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_854_inst_req_1); -- 
    rr_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_858_inst_req_0); -- 
    cr_1700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_858_inst_req_1); -- 
    convTranspose_CP_39_elements(482) <= OrReduce(convTranspose_CP_39_elements(209) & convTranspose_CP_39_elements(122));
    -- CP-element group 483:  transition  output  delay-element  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	221 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	487 
    -- CP-element group 483:  members (5) 
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/$exit
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/$exit
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$exit
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_926_konst_delay_trans
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_req
      -- 
    phi_stmt_920_req_3623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_920_req_3623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(483), ack => phi_stmt_920_req_1); -- 
    -- Element group convTranspose_CP_39_elements(483) is a control-delay.
    cp_element_483_delay: control_delay_element  generic map(name => " 483_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(221), ack => convTranspose_CP_39_elements(483), clk => clk, reset =>reset);
    -- CP-element group 484:  transition  input  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	230 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	486 
    -- CP-element group 484:  members (2) 
      -- CP-element group 484: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/ra
      -- 
    ra_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_0, ack => convTranspose_CP_39_elements(484)); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	230 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	486 
    -- CP-element group 485:  members (2) 
      -- CP-element group 485: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/ca
      -- 
    ca_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_1, ack => convTranspose_CP_39_elements(485)); -- 
    -- CP-element group 486:  join  transition  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	484 
    -- CP-element group 486: 	485 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (6) 
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_req
      -- 
    phi_stmt_920_req_3649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_920_req_3649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(486), ack => phi_stmt_920_req_0); -- 
    convTranspose_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(484) & convTranspose_CP_39_elements(485);
      gj_convTranspose_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  merge  transition  place  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	483 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487:  members (2) 
      -- CP-element group 487: 	 branch_block_stmt_32/merge_stmt_919_PhiReqMerge
      -- CP-element group 487: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(487) <= OrReduce(convTranspose_CP_39_elements(483) & convTranspose_CP_39_elements(486));
    -- CP-element group 488:  fork  transition  place  input  output  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	222 
    -- CP-element group 488: 	223 
    -- CP-element group 488: 	225 
    -- CP-element group 488: 	227 
    -- CP-element group 488:  members (29) 
      -- CP-element group 488: 	 branch_block_stmt_32/merge_stmt_919__exit__
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950__entry__
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_update_start_
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resized_1
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scaled_1
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_computed_1
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/$exit
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/index_resize_req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/index_resize_ack
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/$exit
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/scale_rename_req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/scale_rename_ack
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_update_start
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_update_start_
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/cr
      -- CP-element group 488: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/$exit
      -- CP-element group 488: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/phi_stmt_920_ack
      -- 
    phi_stmt_920_ack_3654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_920_ack_0, ack => convTranspose_CP_39_elements(488)); -- 
    req_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => array_obj_ref_932_index_offset_req_0); -- 
    req_1770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => array_obj_ref_932_index_offset_req_1); -- 
    req_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => addr_of_933_final_reg_req_1); -- 
    cr_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => ptr_deref_936_store_0_req_1); -- 
    -- CP-element group 489:  merge  fork  transition  place  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	219 
    -- CP-element group 489: 	229 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	231 
    -- CP-element group 489: 	232 
    -- CP-element group 489: 	234 
    -- CP-element group 489:  members (16) 
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959__exit__
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968__entry__
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_Sample/crr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/call_stmt_962_Update/ccr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_968/type_cast_967_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959_PhiReqMerge
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/$exit
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/dummy
      -- 
    crr_1866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => call_stmt_962_call_req_0); -- 
    ccr_1871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => call_stmt_962_call_req_1); -- 
    cr_1885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_967_inst_req_1); -- 
    convTranspose_CP_39_elements(489) <= OrReduce(convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(229));
    -- CP-element group 490:  transition  output  delay-element  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	420 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	494 
    -- CP-element group 490:  members (5) 
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/$exit
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1350/$exit
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/$exit
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1354_konst_delay_trans
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_req
      -- 
    phi_stmt_1350_req_3700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1350_req_3700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(490), ack => phi_stmt_1350_req_0); -- 
    -- Element group convTranspose_CP_39_elements(490) is a control-delay.
    cp_element_490_delay: control_delay_element  generic map(name => " 490_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(420), ack => convTranspose_CP_39_elements(490), clk => clk, reset =>reset);
    -- CP-element group 491:  transition  input  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	468 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	493 
    -- CP-element group 491:  members (2) 
      -- CP-element group 491: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/Sample/ra
      -- 
    ra_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_0, ack => convTranspose_CP_39_elements(491)); -- 
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	468 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492:  members (2) 
      -- CP-element group 492: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/Update/ca
      -- 
    ca_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1356_inst_ack_1, ack => convTranspose_CP_39_elements(492)); -- 
    -- CP-element group 493:  join  transition  output  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	491 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (6) 
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_sources/type_cast_1356/SplitProtocol/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1350/phi_stmt_1350_req
      -- 
    phi_stmt_1350_req_3726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1350_req_3726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(493), ack => phi_stmt_1350_req_1); -- 
    convTranspose_cp_element_group_493: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_493"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(491) & convTranspose_CP_39_elements(492);
      gj_convTranspose_cp_element_group_493 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(493), clk => clk, reset => reset); --
    end block;
    -- CP-element group 494:  merge  transition  place  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	490 
    -- CP-element group 494: 	493 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (2) 
      -- CP-element group 494: 	 branch_block_stmt_32/merge_stmt_1349_PhiReqMerge
      -- CP-element group 494: 	 branch_block_stmt_32/merge_stmt_1349_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(494) <= OrReduce(convTranspose_CP_39_elements(490) & convTranspose_CP_39_elements(493));
    -- CP-element group 495:  fork  transition  place  input  output  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	421 
    -- CP-element group 495: 	422 
    -- CP-element group 495: 	424 
    -- CP-element group 495: 	426 
    -- CP-element group 495: 	428 
    -- CP-element group 495: 	430 
    -- CP-element group 495: 	432 
    -- CP-element group 495: 	434 
    -- CP-element group 495: 	436 
    -- CP-element group 495: 	438 
    -- CP-element group 495: 	440 
    -- CP-element group 495: 	442 
    -- CP-element group 495:  members (53) 
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_scale_1/scale_rename_ack
      -- CP-element group 495: 	 branch_block_stmt_32/merge_stmt_1349__exit__
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477__entry__
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_resize_1/index_resize_req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_resize_1/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_resize_1/$exit
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_Sample/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_scale_1/scale_rename_req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_update_start
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_resize_1/index_resize_ack
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_scaled_1
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_computed_1
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_scale_1/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_Update/req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_scale_1/$exit
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_final_index_sum_regn_Sample/req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1371_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/array_obj_ref_1362_index_resized_1
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1431_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1401_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/word_access_complete/word_0/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/word_access_complete/word_0/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/word_access_complete/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1391_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1421_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1441_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/ptr_deref_1367_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_complete/req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1381_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/addr_of_1363_complete/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1364_to_assign_stmt_1477/type_cast_1411_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/merge_stmt_1349_PhiAck/$exit
      -- CP-element group 495: 	 branch_block_stmt_32/merge_stmt_1349_PhiAck/phi_stmt_1350_ack
      -- 
    phi_stmt_1350_ack_3731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1350_ack_0, ack => convTranspose_CP_39_elements(495)); -- 
    cr_3300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1431_inst_req_1); -- 
    req_3137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => array_obj_ref_1362_index_offset_req_1); -- 
    cr_3216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1371_inst_req_1); -- 
    cr_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1401_inst_req_1); -- 
    req_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => array_obj_ref_1362_index_offset_req_0); -- 
    cr_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => ptr_deref_1367_load_0_req_1); -- 
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1391_inst_req_1); -- 
    cr_3314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1441_inst_req_1); -- 
    cr_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1421_inst_req_1); -- 
    cr_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1381_inst_req_1); -- 
    req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => addr_of_1363_final_reg_req_1); -- 
    cr_3272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1411_inst_req_1); -- 
    -- CP-element group 496:  merge  transition  place  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	418 
    -- CP-element group 496: 	467 
    -- CP-element group 496: successors 
    -- CP-element group 496:  members (16) 
      -- CP-element group 496: 	 $exit
      -- CP-element group 496: 	 branch_block_stmt_32/$exit
      -- CP-element group 496: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1486__exit__
      -- CP-element group 496: 	 branch_block_stmt_32/return__
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1488__exit__
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1486_PhiReqMerge
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1486_PhiAck/$entry
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1486_PhiAck/$exit
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1486_PhiAck/dummy
      -- CP-element group 496: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 496: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1488_PhiReqMerge
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1488_PhiAck/$entry
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1488_PhiAck/$exit
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1488_PhiAck/dummy
      -- 
    convTranspose_CP_39_elements(496) <= OrReduce(convTranspose_CP_39_elements(418) & convTranspose_CP_39_elements(467));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar525_931_resized : std_logic_vector(13 downto 0);
    signal R_indvar525_931_scaled : std_logic_vector(13 downto 0);
    signal R_indvar539_687_resized : std_logic_vector(10 downto 0);
    signal R_indvar539_687_scaled : std_logic_vector(10 downto 0);
    signal R_indvar555_480_resized : std_logic_vector(13 downto 0);
    signal R_indvar555_480_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1361_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1361_scaled : std_logic_vector(13 downto 0);
    signal add108_333 : std_logic_vector(15 downto 0);
    signal add117_358 : std_logic_vector(15 downto 0);
    signal add126_383 : std_logic_vector(15 downto 0);
    signal add12_82 : std_logic_vector(15 downto 0);
    signal add135_408 : std_logic_vector(15 downto 0);
    signal add150_508 : std_logic_vector(63 downto 0);
    signal add156_526 : std_logic_vector(63 downto 0);
    signal add162_544 : std_logic_vector(63 downto 0);
    signal add168_562 : std_logic_vector(63 downto 0);
    signal add174_580 : std_logic_vector(63 downto 0);
    signal add180_598 : std_logic_vector(63 downto 0);
    signal add186_616 : std_logic_vector(63 downto 0);
    signal add206_715 : std_logic_vector(63 downto 0);
    signal add212_733 : std_logic_vector(63 downto 0);
    signal add218_751 : std_logic_vector(63 downto 0);
    signal add21_107 : std_logic_vector(15 downto 0);
    signal add224_769 : std_logic_vector(63 downto 0);
    signal add230_787 : std_logic_vector(63 downto 0);
    signal add236_805 : std_logic_vector(63 downto 0);
    signal add242_823 : std_logic_vector(63 downto 0);
    signal add30_132 : std_logic_vector(15 downto 0);
    signal add39_157 : std_logic_vector(15 downto 0);
    signal add48_182 : std_logic_vector(15 downto 0);
    signal add57_207 : std_logic_vector(15 downto 0);
    signal add74_247 : std_logic_vector(31 downto 0);
    signal add79_252 : std_logic_vector(31 downto 0);
    signal add99_308 : std_logic_vector(15 downto 0);
    signal add_57 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1362_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1362_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1362_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1362_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1362_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1362_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_688_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_932_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_690 : std_logic_vector(31 downto 0);
    signal arrayidx269_934 : std_logic_vector(31 downto 0);
    signal arrayidx432_1364 : std_logic_vector(31 downto 0);
    signal arrayidx_483 : std_logic_vector(31 downto 0);
    signal call101_311 : std_logic_vector(7 downto 0);
    signal call106_324 : std_logic_vector(7 downto 0);
    signal call10_73 : std_logic_vector(7 downto 0);
    signal call110_336 : std_logic_vector(7 downto 0);
    signal call115_349 : std_logic_vector(7 downto 0);
    signal call119_361 : std_logic_vector(7 downto 0);
    signal call124_374 : std_logic_vector(7 downto 0);
    signal call128_386 : std_logic_vector(7 downto 0);
    signal call133_399 : std_logic_vector(7 downto 0);
    signal call143_486 : std_logic_vector(7 downto 0);
    signal call147_499 : std_logic_vector(7 downto 0);
    signal call14_85 : std_logic_vector(7 downto 0);
    signal call153_517 : std_logic_vector(7 downto 0);
    signal call159_535 : std_logic_vector(7 downto 0);
    signal call165_553 : std_logic_vector(7 downto 0);
    signal call171_571 : std_logic_vector(7 downto 0);
    signal call177_589 : std_logic_vector(7 downto 0);
    signal call183_607 : std_logic_vector(7 downto 0);
    signal call199_693 : std_logic_vector(7 downto 0);
    signal call19_98 : std_logic_vector(7 downto 0);
    signal call203_706 : std_logic_vector(7 downto 0);
    signal call209_724 : std_logic_vector(7 downto 0);
    signal call215_742 : std_logic_vector(7 downto 0);
    signal call221_760 : std_logic_vector(7 downto 0);
    signal call227_778 : std_logic_vector(7 downto 0);
    signal call233_796 : std_logic_vector(7 downto 0);
    signal call239_814 : std_logic_vector(7 downto 0);
    signal call23_110 : std_logic_vector(7 downto 0);
    signal call275_962 : std_logic_vector(63 downto 0);
    signal call28_123 : std_logic_vector(7 downto 0);
    signal call2_48 : std_logic_vector(7 downto 0);
    signal call32_135 : std_logic_vector(7 downto 0);
    signal call346_1184 : std_logic_vector(15 downto 0);
    signal call348_1187 : std_logic_vector(15 downto 0);
    signal call350_1190 : std_logic_vector(15 downto 0);
    signal call352_1193 : std_logic_vector(15 downto 0);
    signal call354_1196 : std_logic_vector(63 downto 0);
    signal call37_148 : std_logic_vector(7 downto 0);
    signal call41_160 : std_logic_vector(7 downto 0);
    signal call46_173 : std_logic_vector(7 downto 0);
    signal call50_185 : std_logic_vector(7 downto 0);
    signal call55_198 : std_logic_vector(7 downto 0);
    signal call5_60 : std_logic_vector(7 downto 0);
    signal call92_286 : std_logic_vector(7 downto 0);
    signal call97_299 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp194509_430 : std_logic_vector(0 downto 0);
    signal cmp264505_875 : std_logic_vector(0 downto 0);
    signal cmp513_415 : std_logic_vector(0 downto 0);
    signal conv104_315 : std_logic_vector(15 downto 0);
    signal conv107_328 : std_logic_vector(15 downto 0);
    signal conv113_340 : std_logic_vector(15 downto 0);
    signal conv116_353 : std_logic_vector(15 downto 0);
    signal conv11_77 : std_logic_vector(15 downto 0);
    signal conv122_365 : std_logic_vector(15 downto 0);
    signal conv125_378 : std_logic_vector(15 downto 0);
    signal conv131_390 : std_logic_vector(15 downto 0);
    signal conv134_403 : std_logic_vector(15 downto 0);
    signal conv144_490 : std_logic_vector(63 downto 0);
    signal conv149_503 : std_logic_vector(63 downto 0);
    signal conv155_521 : std_logic_vector(63 downto 0);
    signal conv161_539 : std_logic_vector(63 downto 0);
    signal conv167_557 : std_logic_vector(63 downto 0);
    signal conv173_575 : std_logic_vector(63 downto 0);
    signal conv179_593 : std_logic_vector(63 downto 0);
    signal conv17_89 : std_logic_vector(15 downto 0);
    signal conv185_611 : std_logic_vector(63 downto 0);
    signal conv1_39 : std_logic_vector(15 downto 0);
    signal conv200_697 : std_logic_vector(63 downto 0);
    signal conv205_710 : std_logic_vector(63 downto 0);
    signal conv20_102 : std_logic_vector(15 downto 0);
    signal conv211_728 : std_logic_vector(63 downto 0);
    signal conv217_746 : std_logic_vector(63 downto 0);
    signal conv223_764 : std_logic_vector(63 downto 0);
    signal conv229_782 : std_logic_vector(63 downto 0);
    signal conv235_800 : std_logic_vector(63 downto 0);
    signal conv241_818 : std_logic_vector(63 downto 0);
    signal conv253_851 : std_logic_vector(31 downto 0);
    signal conv255_855 : std_logic_vector(31 downto 0);
    signal conv258_859 : std_logic_vector(31 downto 0);
    signal conv26_114 : std_logic_vector(15 downto 0);
    signal conv276_968 : std_logic_vector(63 downto 0);
    signal conv29_127 : std_logic_vector(15 downto 0);
    signal conv305_1050 : std_logic_vector(15 downto 0);
    signal conv307_1057 : std_logic_vector(15 downto 0);
    signal conv322_1106 : std_logic_vector(15 downto 0);
    signal conv324_1113 : std_logic_vector(15 downto 0);
    signal conv339_1162 : std_logic_vector(15 downto 0);
    signal conv341_1169 : std_logic_vector(15 downto 0);
    signal conv355_1201 : std_logic_vector(63 downto 0);
    signal conv35_139 : std_logic_vector(15 downto 0);
    signal conv361_1210 : std_logic_vector(7 downto 0);
    signal conv367_1220 : std_logic_vector(7 downto 0);
    signal conv373_1230 : std_logic_vector(7 downto 0);
    signal conv379_1240 : std_logic_vector(7 downto 0);
    signal conv385_1250 : std_logic_vector(7 downto 0);
    signal conv38_152 : std_logic_vector(15 downto 0);
    signal conv391_1260 : std_logic_vector(7 downto 0);
    signal conv397_1270 : std_logic_vector(7 downto 0);
    signal conv3_52 : std_logic_vector(15 downto 0);
    signal conv403_1280 : std_logic_vector(7 downto 0);
    signal conv437_1372 : std_logic_vector(7 downto 0);
    signal conv443_1382 : std_logic_vector(7 downto 0);
    signal conv449_1392 : std_logic_vector(7 downto 0);
    signal conv44_164 : std_logic_vector(15 downto 0);
    signal conv455_1402 : std_logic_vector(7 downto 0);
    signal conv461_1412 : std_logic_vector(7 downto 0);
    signal conv467_1422 : std_logic_vector(7 downto 0);
    signal conv473_1432 : std_logic_vector(7 downto 0);
    signal conv479_1442 : std_logic_vector(7 downto 0);
    signal conv47_177 : std_logic_vector(15 downto 0);
    signal conv53_189 : std_logic_vector(15 downto 0);
    signal conv56_202 : std_logic_vector(15 downto 0);
    signal conv61_211 : std_logic_vector(31 downto 0);
    signal conv63_215 : std_logic_vector(31 downto 0);
    signal conv65_219 : std_logic_vector(31 downto 0);
    signal conv82_256 : std_logic_vector(31 downto 0);
    signal conv84_260 : std_logic_vector(31 downto 0);
    signal conv87_264 : std_logic_vector(31 downto 0);
    signal conv8_64 : std_logic_vector(15 downto 0);
    signal conv90_268 : std_logic_vector(31 downto 0);
    signal conv95_290 : std_logic_vector(15 downto 0);
    signal conv98_303 : std_logic_vector(15 downto 0);
    signal exitcond1_1477 : std_logic_vector(0 downto 0);
    signal exitcond2_838 : std_logic_vector(0 downto 0);
    signal exitcond3_631 : std_logic_vector(0 downto 0);
    signal exitcond_950 : std_logic_vector(0 downto 0);
    signal iNsTr_14_241 : std_logic_vector(31 downto 0);
    signal iNsTr_195_1334 : std_logic_vector(63 downto 0);
    signal iNsTr_26_453 : std_logic_vector(63 downto 0);
    signal iNsTr_39_660 : std_logic_vector(63 downto 0);
    signal iNsTr_53_904 : std_logic_vector(63 downto 0);
    signal indvar525_920 : std_logic_vector(63 downto 0);
    signal indvar539_676 : std_logic_vector(63 downto 0);
    signal indvar555_469 : std_logic_vector(63 downto 0);
    signal indvar_1350 : std_logic_vector(63 downto 0);
    signal indvarx_xnext526_945 : std_logic_vector(63 downto 0);
    signal indvarx_xnext540_833 : std_logic_vector(63 downto 0);
    signal indvarx_xnext556_626 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1472 : std_logic_vector(63 downto 0);
    signal mul256_864 : std_logic_vector(31 downto 0);
    signal mul259_869 : std_logic_vector(31 downto 0);
    signal mul66_229 : std_logic_vector(31 downto 0);
    signal mul85_273 : std_logic_vector(31 downto 0);
    signal mul88_278 : std_logic_vector(31 downto 0);
    signal mul91_283 : std_logic_vector(31 downto 0);
    signal mul_224 : std_logic_vector(31 downto 0);
    signal ptr_deref_1367_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1367_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1367_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1367_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1367_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_618_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_618_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_618_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_618_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_618_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_618_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_825_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_825_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_825_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_825_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_825_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_825_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_936_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_936_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_936_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_936_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_936_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_936_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_321 : std_logic_vector(15 downto 0);
    signal shl114_346 : std_logic_vector(15 downto 0);
    signal shl123_371 : std_logic_vector(15 downto 0);
    signal shl132_396 : std_logic_vector(15 downto 0);
    signal shl146_496 : std_logic_vector(63 downto 0);
    signal shl152_514 : std_logic_vector(63 downto 0);
    signal shl158_532 : std_logic_vector(63 downto 0);
    signal shl164_550 : std_logic_vector(63 downto 0);
    signal shl170_568 : std_logic_vector(63 downto 0);
    signal shl176_586 : std_logic_vector(63 downto 0);
    signal shl182_604 : std_logic_vector(63 downto 0);
    signal shl18_95 : std_logic_vector(15 downto 0);
    signal shl202_703 : std_logic_vector(63 downto 0);
    signal shl208_721 : std_logic_vector(63 downto 0);
    signal shl214_739 : std_logic_vector(63 downto 0);
    signal shl220_757 : std_logic_vector(63 downto 0);
    signal shl226_775 : std_logic_vector(63 downto 0);
    signal shl232_793 : std_logic_vector(63 downto 0);
    signal shl238_811 : std_logic_vector(63 downto 0);
    signal shl27_120 : std_logic_vector(15 downto 0);
    signal shl36_145 : std_logic_vector(15 downto 0);
    signal shl45_170 : std_logic_vector(15 downto 0);
    signal shl54_195 : std_logic_vector(15 downto 0);
    signal shl96_296 : std_logic_vector(15 downto 0);
    signal shl9_70 : std_logic_vector(15 downto 0);
    signal shl_45 : std_logic_vector(15 downto 0);
    signal shr304_1046 : std_logic_vector(31 downto 0);
    signal shr321_1102 : std_logic_vector(31 downto 0);
    signal shr338_1158 : std_logic_vector(31 downto 0);
    signal shr364_1216 : std_logic_vector(63 downto 0);
    signal shr370_1226 : std_logic_vector(63 downto 0);
    signal shr376_1236 : std_logic_vector(63 downto 0);
    signal shr382_1246 : std_logic_vector(63 downto 0);
    signal shr388_1256 : std_logic_vector(63 downto 0);
    signal shr394_1266 : std_logic_vector(63 downto 0);
    signal shr400_1276 : std_logic_vector(63 downto 0);
    signal shr440_1378 : std_logic_vector(63 downto 0);
    signal shr446_1388 : std_logic_vector(63 downto 0);
    signal shr452_1398 : std_logic_vector(63 downto 0);
    signal shr458_1408 : std_logic_vector(63 downto 0);
    signal shr464_1418 : std_logic_vector(63 downto 0);
    signal shr470_1428 : std_logic_vector(63 downto 0);
    signal shr476_1438 : std_logic_vector(63 downto 0);
    signal shr_235 : std_logic_vector(31 downto 0);
    signal sub_1206 : std_logic_vector(63 downto 0);
    signal tmp433_1368 : std_logic_vector(63 downto 0);
    signal tmp520_1318 : std_logic_vector(31 downto 0);
    signal tmp520x_xop_1330 : std_logic_vector(31 downto 0);
    signal tmp521_1324 : std_logic_vector(0 downto 0);
    signal tmp524_1347 : std_logic_vector(63 downto 0);
    signal tmp532_888 : std_logic_vector(31 downto 0);
    signal tmp532x_xop_900 : std_logic_vector(31 downto 0);
    signal tmp533_894 : std_logic_vector(0 downto 0);
    signal tmp537_917 : std_logic_vector(63 downto 0);
    signal tmp548_644 : std_logic_vector(31 downto 0);
    signal tmp548x_xop_656 : std_logic_vector(31 downto 0);
    signal tmp549_650 : std_logic_vector(0 downto 0);
    signal tmp553_673 : std_logic_vector(63 downto 0);
    signal tmp562x_xop_449 : std_logic_vector(31 downto 0);
    signal tmp563_443 : std_logic_vector(0 downto 0);
    signal tmp567_466 : std_logic_vector(63 downto 0);
    signal type_cast_1003_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1044_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1100_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1156_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1199_wire : std_logic_vector(63 downto 0);
    signal type_cast_1214_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1224_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1234_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1244_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1264_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1274_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1316_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1322_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1328_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1345_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1354_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1356_wire : std_logic_vector(63 downto 0);
    signal type_cast_1376_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1386_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1396_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1406_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1416_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1426_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1436_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_143_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1470_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_168_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_193_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_245_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_294_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_319_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_344_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_369_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_394_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_412_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_428_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_43_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_441_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_447_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_464_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_473_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_475_wire : std_logic_vector(63 downto 0);
    signal type_cast_494_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_530_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_548_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_584_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_602_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_642_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_664_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_671_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_679_wire : std_logic_vector(63 downto 0);
    signal type_cast_682_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_701_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_719_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_737_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_791_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_809_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_831_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_873_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_898_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_915_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_923_wire : std_logic_vector(63 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_938_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_93_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_966_wire : std_logic_vector(63 downto 0);
    signal type_cast_999_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop569_910 : std_logic_vector(63 downto 0);
    signal xx_xop570_666 : std_logic_vector(63 downto 0);
    signal xx_xop571_459 : std_logic_vector(63 downto 0);
    signal xx_xop_1340 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1362_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1362_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1362_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1362_resized_base_address <= "00000000000000";
    array_obj_ref_481_constant_part_of_offset <= "00000000000000";
    array_obj_ref_481_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_481_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_481_resized_base_address <= "00000000000000";
    array_obj_ref_688_constant_part_of_offset <= "00000100010";
    array_obj_ref_688_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_688_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_688_resized_base_address <= "00000000000";
    array_obj_ref_932_constant_part_of_offset <= "00000000000000";
    array_obj_ref_932_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_932_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_932_resized_base_address <= "00000000000000";
    ptr_deref_1367_word_offset_0 <= "00000000000000";
    ptr_deref_618_word_offset_0 <= "00000000000000";
    ptr_deref_825_word_offset_0 <= "00000000000";
    ptr_deref_936_word_offset_0 <= "00000000000000";
    type_cast_1003_wire_constant <= "0000000000000000";
    type_cast_1044_wire_constant <= "00000000000000000000000000010010";
    type_cast_1100_wire_constant <= "00000000000000000000000000010001";
    type_cast_1156_wire_constant <= "00000000000000000000000000010000";
    type_cast_118_wire_constant <= "0000000000001000";
    type_cast_1214_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1224_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1234_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1244_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1254_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1264_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1274_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1316_wire_constant <= "00000000000000000000000000000010";
    type_cast_1322_wire_constant <= "00000000000000000000000000000001";
    type_cast_1328_wire_constant <= "11111111111111111111111111111111";
    type_cast_1338_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1345_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1354_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1376_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1396_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1406_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1416_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1426_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1436_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_143_wire_constant <= "0000000000001000";
    type_cast_1470_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_168_wire_constant <= "0000000000001000";
    type_cast_193_wire_constant <= "0000000000001000";
    type_cast_233_wire_constant <= "00000000000000000000000000000010";
    type_cast_239_wire_constant <= "00000000000000000000000000000001";
    type_cast_245_wire_constant <= "01111111111111111111111111111110";
    type_cast_294_wire_constant <= "0000000000001000";
    type_cast_319_wire_constant <= "0000000000001000";
    type_cast_344_wire_constant <= "0000000000001000";
    type_cast_369_wire_constant <= "0000000000001000";
    type_cast_394_wire_constant <= "0000000000001000";
    type_cast_412_wire_constant <= "00000000000000000000000000000011";
    type_cast_428_wire_constant <= "00000000000000000000000000000011";
    type_cast_43_wire_constant <= "0000000000001000";
    type_cast_441_wire_constant <= "00000000000000000000000000000001";
    type_cast_447_wire_constant <= "11111111111111111111111111111111";
    type_cast_457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_464_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_473_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_494_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_512_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_530_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_548_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_566_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_584_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_602_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_624_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_642_wire_constant <= "00000000000000000000000000000010";
    type_cast_648_wire_constant <= "00000000000000000000000000000001";
    type_cast_654_wire_constant <= "11111111111111111111111111111111";
    type_cast_664_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_671_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_682_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_68_wire_constant <= "0000000000001000";
    type_cast_701_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_719_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_737_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_791_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_809_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_831_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_873_wire_constant <= "00000000000000000000000000000011";
    type_cast_886_wire_constant <= "00000000000000000000000000000010";
    type_cast_892_wire_constant <= "00000000000000000000000000000001";
    type_cast_898_wire_constant <= "11111111111111111111111111111111";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_915_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_926_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_938_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_93_wire_constant <= "0000000000001000";
    type_cast_943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_999_wire_constant <= "0000000000000000";
    phi_stmt_1350: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1354_wire_constant & type_cast_1356_wire;
      req <= phi_stmt_1350_req_0 & phi_stmt_1350_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1350",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1350_ack_0,
          idata => idata,
          odata => indvar_1350,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1350
    phi_stmt_469: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_473_wire_constant & type_cast_475_wire;
      req <= phi_stmt_469_req_0 & phi_stmt_469_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_469",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_469_ack_0,
          idata => idata,
          odata => indvar555_469,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_469
    phi_stmt_676: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_679_wire & type_cast_682_wire_constant;
      req <= phi_stmt_676_req_0 & phi_stmt_676_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_676",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_676_ack_0,
          idata => idata,
          odata => indvar539_676,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_676
    phi_stmt_920: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_923_wire & type_cast_926_wire_constant;
      req <= phi_stmt_920_req_0 & phi_stmt_920_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_920",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_920_ack_0,
          idata => idata,
          odata => indvar525_920,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_920
    -- flow-through select operator MUX_1346_inst
    tmp524_1347 <= xx_xop_1340 when (tmp521_1324(0) /=  '0') else type_cast_1345_wire_constant;
    -- flow-through select operator MUX_465_inst
    tmp567_466 <= xx_xop571_459 when (tmp563_443(0) /=  '0') else type_cast_464_wire_constant;
    -- flow-through select operator MUX_672_inst
    tmp553_673 <= xx_xop570_666 when (tmp549_650(0) /=  '0') else type_cast_671_wire_constant;
    -- flow-through select operator MUX_916_inst
    tmp537_917 <= xx_xop569_910 when (tmp533_894(0) /=  '0') else type_cast_915_wire_constant;
    addr_of_1363_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1363_final_reg_req_0;
      addr_of_1363_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1363_final_reg_req_1;
      addr_of_1363_final_reg_ack_1<= rack(0);
      addr_of_1363_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1363_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1362_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx432_1364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_482_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_482_final_reg_req_0;
      addr_of_482_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_482_final_reg_req_1;
      addr_of_482_final_reg_ack_1<= rack(0);
      addr_of_482_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_482_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_481_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_689_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_689_final_reg_req_0;
      addr_of_689_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_689_final_reg_req_1;
      addr_of_689_final_reg_ack_1<= rack(0);
      addr_of_689_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_689_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_688_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_933_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_933_final_reg_req_0;
      addr_of_933_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_933_final_reg_req_1;
      addr_of_933_final_reg_ack_1<= rack(0);
      addr_of_933_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_933_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_932_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_101_inst_req_0;
      type_cast_101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_101_inst_req_1;
      type_cast_101_inst_ack_1<= rack(0);
      type_cast_101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1049_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1049_inst_req_0;
      type_cast_1049_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1049_inst_req_1;
      type_cast_1049_inst_ack_1<= rack(0);
      type_cast_1049_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1049_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1046,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1050,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1056_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1056_inst_req_0;
      type_cast_1056_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1056_inst_req_1;
      type_cast_1056_inst_ack_1<= rack(0);
      type_cast_1056_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1056_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1105_inst_req_0;
      type_cast_1105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1105_inst_req_1;
      type_cast_1105_inst_ack_1<= rack(0);
      type_cast_1105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr321_1102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1112_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1112_inst_req_0;
      type_cast_1112_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1112_inst_req_1;
      type_cast_1112_inst_ack_1<= rack(0);
      type_cast_1112_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1112_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1113,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1161_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1161_inst_req_0;
      type_cast_1161_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1161_inst_req_1;
      type_cast_1161_inst_ack_1<= rack(0);
      type_cast_1161_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1161_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1162,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1168_inst_req_0;
      type_cast_1168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1168_inst_req_1;
      type_cast_1168_inst_ack_1<= rack(0);
      type_cast_1168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1200_inst_req_0;
      type_cast_1200_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1200_inst_req_1;
      type_cast_1200_inst_ack_1<= rack(0);
      type_cast_1200_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1200_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1199_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1209_inst_req_0;
      type_cast_1209_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1209_inst_req_1;
      type_cast_1209_inst_ack_1<= rack(0);
      type_cast_1209_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1209_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1206,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv361_1210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1219_inst_req_0;
      type_cast_1219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1219_inst_req_1;
      type_cast_1219_inst_ack_1<= rack(0);
      type_cast_1219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr364_1216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv367_1220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1229_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1229_inst_req_0;
      type_cast_1229_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1229_inst_req_1;
      type_cast_1229_inst_ack_1<= rack(0);
      type_cast_1229_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1229_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr370_1226,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv373_1230,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1239_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1239_inst_req_0;
      type_cast_1239_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1239_inst_req_1;
      type_cast_1239_inst_ack_1<= rack(0);
      type_cast_1239_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1239_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr376_1236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv379_1240,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1249_inst_req_0;
      type_cast_1249_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1249_inst_req_1;
      type_cast_1249_inst_ack_1<= rack(0);
      type_cast_1249_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1249_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr382_1246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv385_1250,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1259_inst_req_0;
      type_cast_1259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1259_inst_req_1;
      type_cast_1259_inst_ack_1<= rack(0);
      type_cast_1259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr388_1256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv391_1260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1269_inst_req_0;
      type_cast_1269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1269_inst_req_1;
      type_cast_1269_inst_ack_1<= rack(0);
      type_cast_1269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr394_1266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv397_1270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1279_inst_req_0;
      type_cast_1279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1279_inst_req_1;
      type_cast_1279_inst_ack_1<= rack(0);
      type_cast_1279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr400_1276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv403_1280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1333_inst_req_0;
      type_cast_1333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1333_inst_req_1;
      type_cast_1333_inst_ack_1<= rack(0);
      type_cast_1333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp520x_xop_1330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_195_1334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1356_inst_req_0;
      type_cast_1356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1356_inst_req_1;
      type_cast_1356_inst_ack_1<= rack(0);
      type_cast_1356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1472,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1356_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1371_inst_req_0;
      type_cast_1371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1371_inst_req_1;
      type_cast_1371_inst_ack_1<= rack(0);
      type_cast_1371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp433_1368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv437_1372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1381_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1381_inst_req_0;
      type_cast_1381_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1381_inst_req_1;
      type_cast_1381_inst_ack_1<= rack(0);
      type_cast_1381_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1381_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr440_1378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv443_1382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_138_inst_req_0;
      type_cast_138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_138_inst_req_1;
      type_cast_138_inst_ack_1<= rack(0);
      type_cast_138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1391_inst_req_0;
      type_cast_1391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1391_inst_req_1;
      type_cast_1391_inst_ack_1<= rack(0);
      type_cast_1391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr446_1388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv449_1392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1401_inst_req_0;
      type_cast_1401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1401_inst_req_1;
      type_cast_1401_inst_ack_1<= rack(0);
      type_cast_1401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr452_1398,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv455_1402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1411_inst_req_0;
      type_cast_1411_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1411_inst_req_1;
      type_cast_1411_inst_ack_1<= rack(0);
      type_cast_1411_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1411_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr458_1408,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv461_1412,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1421_inst_req_0;
      type_cast_1421_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1421_inst_req_1;
      type_cast_1421_inst_ack_1<= rack(0);
      type_cast_1421_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1421_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr464_1418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv467_1422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1431_inst_req_0;
      type_cast_1431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1431_inst_req_1;
      type_cast_1431_inst_ack_1<= rack(0);
      type_cast_1431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr470_1428,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv473_1432,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1441_inst_req_0;
      type_cast_1441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1441_inst_req_1;
      type_cast_1441_inst_ack_1<= rack(0);
      type_cast_1441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr476_1438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv479_1442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_151_inst_req_0;
      type_cast_151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_151_inst_req_1;
      type_cast_151_inst_ack_1<= rack(0);
      type_cast_151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_163_inst_req_0;
      type_cast_163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_163_inst_req_1;
      type_cast_163_inst_ack_1<= rack(0);
      type_cast_163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_176_inst_req_0;
      type_cast_176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_176_inst_req_1;
      type_cast_176_inst_ack_1<= rack(0);
      type_cast_176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_188_inst_req_0;
      type_cast_188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_188_inst_req_1;
      type_cast_188_inst_ack_1<= rack(0);
      type_cast_188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_201_inst_req_0;
      type_cast_201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_201_inst_req_1;
      type_cast_201_inst_ack_1<= rack(0);
      type_cast_201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_210_inst_req_0;
      type_cast_210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_210_inst_req_1;
      type_cast_210_inst_ack_1<= rack(0);
      type_cast_210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_57,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_214_inst_req_0;
      type_cast_214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_214_inst_req_1;
      type_cast_214_inst_ack_1<= rack(0);
      type_cast_214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_82,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_218_inst_req_0;
      type_cast_218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_218_inst_req_1;
      type_cast_218_inst_ack_1<= rack(0);
      type_cast_218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_255_inst_req_0;
      type_cast_255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_255_inst_req_1;
      type_cast_255_inst_ack_1<= rack(0);
      type_cast_255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_259_inst_req_0;
      type_cast_259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_259_inst_req_1;
      type_cast_259_inst_ack_1<= rack(0);
      type_cast_259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_263_inst_req_0;
      type_cast_263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_263_inst_req_1;
      type_cast_263_inst_ack_1<= rack(0);
      type_cast_263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_267_inst_req_0;
      type_cast_267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_267_inst_req_1;
      type_cast_267_inst_ack_1<= rack(0);
      type_cast_267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_268,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_289_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_289_inst_req_0;
      type_cast_289_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_289_inst_req_1;
      type_cast_289_inst_ack_1<= rack(0);
      type_cast_289_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_289_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_290,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_302_inst_req_0;
      type_cast_302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_302_inst_req_1;
      type_cast_302_inst_ack_1<= rack(0);
      type_cast_302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_314_inst_req_0;
      type_cast_314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_314_inst_req_1;
      type_cast_314_inst_ack_1<= rack(0);
      type_cast_314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_327_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_327_inst_req_0;
      type_cast_327_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_327_inst_req_1;
      type_cast_327_inst_ack_1<= rack(0);
      type_cast_327_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_327_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_324,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_328,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_339_inst_req_0;
      type_cast_339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_339_inst_req_1;
      type_cast_339_inst_ack_1<= rack(0);
      type_cast_339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_352_inst_req_0;
      type_cast_352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_352_inst_req_1;
      type_cast_352_inst_ack_1<= rack(0);
      type_cast_352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_364_inst_req_0;
      type_cast_364_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_364_inst_req_1;
      type_cast_364_inst_ack_1<= rack(0);
      type_cast_364_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_364_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_361,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_377_inst_req_0;
      type_cast_377_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_377_inst_req_1;
      type_cast_377_inst_ack_1<= rack(0);
      type_cast_377_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_378,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_389_inst_req_0;
      type_cast_389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_389_inst_req_1;
      type_cast_389_inst_ack_1<= rack(0);
      type_cast_389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_402_inst_req_0;
      type_cast_402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_402_inst_req_1;
      type_cast_402_inst_ack_1<= rack(0);
      type_cast_402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_399,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_452_inst_req_0;
      type_cast_452_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_452_inst_req_1;
      type_cast_452_inst_ack_1<= rack(0);
      type_cast_452_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp562x_xop_449,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_475_inst_req_0;
      type_cast_475_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_475_inst_req_1;
      type_cast_475_inst_ack_1<= rack(0);
      type_cast_475_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext556_626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_475_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_489_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_489_inst_req_0;
      type_cast_489_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_489_inst_req_1;
      type_cast_489_inst_ack_1<= rack(0);
      type_cast_489_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_489_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_486,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_502_inst_req_0;
      type_cast_502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_502_inst_req_1;
      type_cast_502_inst_ack_1<= rack(0);
      type_cast_502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_51_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_51_inst_req_0;
      type_cast_51_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_51_inst_req_1;
      type_cast_51_inst_ack_1<= rack(0);
      type_cast_51_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_51_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_48,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_52,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_520_inst_req_0;
      type_cast_520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_520_inst_req_1;
      type_cast_520_inst_ack_1<= rack(0);
      type_cast_520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_538_inst_req_0;
      type_cast_538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_538_inst_req_1;
      type_cast_538_inst_ack_1<= rack(0);
      type_cast_538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_556_inst_req_0;
      type_cast_556_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_556_inst_req_1;
      type_cast_556_inst_ack_1<= rack(0);
      type_cast_556_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_556_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_557,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_574_inst_req_0;
      type_cast_574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_574_inst_req_1;
      type_cast_574_inst_ack_1<= rack(0);
      type_cast_574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_592_inst_req_0;
      type_cast_592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_592_inst_req_1;
      type_cast_592_inst_ack_1<= rack(0);
      type_cast_592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_610_inst_req_0;
      type_cast_610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_610_inst_req_1;
      type_cast_610_inst_ack_1<= rack(0);
      type_cast_610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_659_inst_req_0;
      type_cast_659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_659_inst_req_1;
      type_cast_659_inst_ack_1<= rack(0);
      type_cast_659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp548x_xop_656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_660,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_679_inst_req_0;
      type_cast_679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_679_inst_req_1;
      type_cast_679_inst_ack_1<= rack(0);
      type_cast_679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext540_833,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_679_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_696_inst_req_0;
      type_cast_696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_696_inst_req_1;
      type_cast_696_inst_ack_1<= rack(0);
      type_cast_696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_693,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_697,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_709_inst_req_0;
      type_cast_709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_709_inst_req_1;
      type_cast_709_inst_ack_1<= rack(0);
      type_cast_709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1<= rack(0);
      type_cast_727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_745_inst_req_0;
      type_cast_745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_745_inst_req_1;
      type_cast_745_inst_ack_1<= rack(0);
      type_cast_745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_742,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_746,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_763_inst_req_0;
      type_cast_763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_763_inst_req_1;
      type_cast_763_inst_ack_1<= rack(0);
      type_cast_763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_760,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_781_inst_req_0;
      type_cast_781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_781_inst_req_1;
      type_cast_781_inst_ack_1<= rack(0);
      type_cast_781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_799_inst_req_0;
      type_cast_799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_799_inst_req_1;
      type_cast_799_inst_ack_1<= rack(0);
      type_cast_799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_800,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_817_inst_req_0;
      type_cast_817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_817_inst_req_1;
      type_cast_817_inst_ack_1<= rack(0);
      type_cast_817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_850_inst_req_0;
      type_cast_850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_850_inst_req_1;
      type_cast_850_inst_ack_1<= rack(0);
      type_cast_850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_854_inst_req_1;
      type_cast_854_inst_ack_1<= rack(0);
      type_cast_854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_858_inst_req_0;
      type_cast_858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_858_inst_req_1;
      type_cast_858_inst_ack_1<= rack(0);
      type_cast_858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_408,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_903_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_903_inst_req_0;
      type_cast_903_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_903_inst_req_1;
      type_cast_903_inst_ack_1<= rack(0);
      type_cast_903_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_903_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp532x_xop_900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_923_inst_req_0;
      type_cast_923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_923_inst_req_1;
      type_cast_923_inst_ack_1<= rack(0);
      type_cast_923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext526_945,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_967_inst_req_0;
      type_cast_967_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_967_inst_req_1;
      type_cast_967_inst_ack_1<= rack(0);
      type_cast_967_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_967_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_966_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1362_index_1_rename
    process(R_indvar_1361_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1361_resized;
      ov(13 downto 0) := iv;
      R_indvar_1361_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1362_index_1_resize
    process(indvar_1350) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1350;
      ov := iv(13 downto 0);
      R_indvar_1361_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1362_root_address_inst
    process(array_obj_ref_1362_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1362_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1362_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_index_1_rename
    process(R_indvar555_480_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar555_480_resized;
      ov(13 downto 0) := iv;
      R_indvar555_480_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_index_1_resize
    process(indvar555_469) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar555_469;
      ov := iv(13 downto 0);
      R_indvar555_480_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_root_address_inst
    process(array_obj_ref_481_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_481_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_481_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_index_1_rename
    process(R_indvar539_687_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar539_687_resized;
      ov(10 downto 0) := iv;
      R_indvar539_687_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_index_1_resize
    process(indvar539_676) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar539_676;
      ov := iv(10 downto 0);
      R_indvar539_687_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_root_address_inst
    process(array_obj_ref_688_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_688_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_688_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_index_1_rename
    process(R_indvar525_931_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar525_931_resized;
      ov(13 downto 0) := iv;
      R_indvar525_931_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_index_1_resize
    process(indvar525_920) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar525_920;
      ov := iv(13 downto 0);
      R_indvar525_931_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_root_address_inst
    process(array_obj_ref_932_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_932_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_932_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1367_addr_0
    process(ptr_deref_1367_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1367_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1367_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1367_base_resize
    process(arrayidx432_1364) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx432_1364;
      ov := iv(13 downto 0);
      ptr_deref_1367_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1367_gather_scatter
    process(ptr_deref_1367_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1367_data_0;
      ov(63 downto 0) := iv;
      tmp433_1368 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1367_root_address_inst
    process(ptr_deref_1367_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1367_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1367_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_addr_0
    process(ptr_deref_618_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_618_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_618_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_base_resize
    process(arrayidx_483) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_483;
      ov := iv(13 downto 0);
      ptr_deref_618_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_gather_scatter
    process(add186_616) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_616;
      ov(63 downto 0) := iv;
      ptr_deref_618_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_root_address_inst
    process(ptr_deref_618_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_618_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_618_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_addr_0
    process(ptr_deref_825_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_825_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_825_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_base_resize
    process(arrayidx246_690) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_690;
      ov := iv(10 downto 0);
      ptr_deref_825_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_gather_scatter
    process(add242_823) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_823;
      ov(63 downto 0) := iv;
      ptr_deref_825_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_root_address_inst
    process(ptr_deref_825_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_825_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_825_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_addr_0
    process(ptr_deref_936_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_936_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_base_resize
    process(arrayidx269_934) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_934;
      ov := iv(13 downto 0);
      ptr_deref_936_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_gather_scatter
    process(type_cast_938_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_938_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_936_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_root_address_inst
    process(ptr_deref_936_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_936_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1306_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_875;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1306_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1306_branch_req_0,
          ack0 => if_stmt_1306_branch_ack_0,
          ack1 => if_stmt_1306_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1478_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1477;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1478_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1478_branch_req_0,
          ack0 => if_stmt_1478_branch_ack_0,
          ack1 => if_stmt_1478_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_416_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp513_415;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_416_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_416_branch_req_0,
          ack0 => if_stmt_416_branch_ack_0,
          ack1 => if_stmt_416_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_431_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194509_430;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_431_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_431_branch_req_0,
          ack0 => if_stmt_431_branch_ack_0,
          ack1 => if_stmt_431_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_632_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_631;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_632_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_632_branch_req_0,
          ack0 => if_stmt_632_branch_ack_0,
          ack1 => if_stmt_632_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_839_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_838;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_839_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_839_branch_req_0,
          ack0 => if_stmt_839_branch_ack_0,
          ack1 => if_stmt_839_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_876_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_875;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_876_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_876_branch_req_0,
          ack0 => if_stmt_876_branch_ack_0,
          ack1 => if_stmt_876_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_951_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_950;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_951_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_951_branch_req_0,
          ack0 => if_stmt_951_branch_ack_0,
          ack1 => if_stmt_951_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1329_inst
    process(tmp520_1318) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp520_1318, type_cast_1328_wire_constant, tmp_var);
      tmp520x_xop_1330 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_251_inst
    process(add74_247, shr_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_247, shr_235, tmp_var);
      add79_252 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_448_inst
    process(shr_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_235, type_cast_447_wire_constant, tmp_var);
      tmp562x_xop_449 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_655_inst
    process(tmp548_644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp548_644, type_cast_654_wire_constant, tmp_var);
      tmp548x_xop_656 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_899_inst
    process(tmp532_888) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp532_888, type_cast_898_wire_constant, tmp_var);
      tmp532x_xop_900 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1339_inst
    process(iNsTr_195_1334) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_195_1334, type_cast_1338_wire_constant, tmp_var);
      xx_xop_1340 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1471_inst
    process(indvar_1350) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1350, type_cast_1470_wire_constant, tmp_var);
      indvarx_xnext_1472 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_458_inst
    process(iNsTr_26_453) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_453, type_cast_457_wire_constant, tmp_var);
      xx_xop571_459 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_625_inst
    process(indvar555_469) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar555_469, type_cast_624_wire_constant, tmp_var);
      indvarx_xnext556_626 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_665_inst
    process(iNsTr_39_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_660, type_cast_664_wire_constant, tmp_var);
      xx_xop570_666 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_832_inst
    process(indvar539_676) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar539_676, type_cast_831_wire_constant, tmp_var);
      indvarx_xnext540_833 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_909_inst
    process(iNsTr_53_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_904, type_cast_908_wire_constant, tmp_var);
      xx_xop569_910 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_944_inst
    process(indvar525_920) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar525_920, type_cast_943_wire_constant, tmp_var);
      indvarx_xnext526_945 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_246_inst
    process(iNsTr_14_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_241, type_cast_245_wire_constant, tmp_var);
      add74_247 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1476_inst
    process(indvarx_xnext_1472, tmp524_1347) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1472, tmp524_1347, tmp_var);
      exitcond1_1477 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_630_inst
    process(indvarx_xnext556_626, tmp567_466) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext556_626, tmp567_466, tmp_var);
      exitcond3_631 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_837_inst
    process(indvarx_xnext540_833, tmp553_673) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext540_833, tmp553_673, tmp_var);
      exitcond2_838 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_949_inst
    process(indvarx_xnext526_945, tmp537_917) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext526_945, tmp537_917, tmp_var);
      exitcond_950 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1045_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_1044_wire_constant, tmp_var);
      shr304_1046 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1101_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_1100_wire_constant, tmp_var);
      shr321_1102 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1157_inst
    process(add79_252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_252, type_cast_1156_wire_constant, tmp_var);
      shr338_1158 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1317_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_869, type_cast_1316_wire_constant, tmp_var);
      tmp520_1318 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_234_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_233_wire_constant, tmp_var);
      shr_235 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_240_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_239_wire_constant, tmp_var);
      iNsTr_14_241 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_643_inst
    process(mul91_283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_283, type_cast_642_wire_constant, tmp_var);
      tmp548_644 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_887_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_869, type_cast_886_wire_constant, tmp_var);
      tmp532_888 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1215_inst
    process(sub_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1206, type_cast_1214_wire_constant, tmp_var);
      shr364_1216 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1225_inst
    process(sub_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1206, type_cast_1224_wire_constant, tmp_var);
      shr370_1226 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1235_inst
    process(sub_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1206, type_cast_1234_wire_constant, tmp_var);
      shr376_1236 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1245_inst
    process(sub_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1206, type_cast_1244_wire_constant, tmp_var);
      shr382_1246 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1255_inst
    process(sub_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1206, type_cast_1254_wire_constant, tmp_var);
      shr388_1256 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1265_inst
    process(sub_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1206, type_cast_1264_wire_constant, tmp_var);
      shr394_1266 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1275_inst
    process(sub_1206) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1206, type_cast_1274_wire_constant, tmp_var);
      shr400_1276 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1377_inst
    process(tmp433_1368) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1368, type_cast_1376_wire_constant, tmp_var);
      shr440_1378 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1387_inst
    process(tmp433_1368) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1368, type_cast_1386_wire_constant, tmp_var);
      shr446_1388 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1397_inst
    process(tmp433_1368) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1368, type_cast_1396_wire_constant, tmp_var);
      shr452_1398 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1407_inst
    process(tmp433_1368) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1368, type_cast_1406_wire_constant, tmp_var);
      shr458_1408 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1417_inst
    process(tmp433_1368) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1368, type_cast_1416_wire_constant, tmp_var);
      shr464_1418 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1427_inst
    process(tmp433_1368) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1368, type_cast_1426_wire_constant, tmp_var);
      shr470_1428 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1437_inst
    process(tmp433_1368) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1368, type_cast_1436_wire_constant, tmp_var);
      shr476_1438 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_223_inst
    process(conv63_215, conv61_211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_215, conv61_211, tmp_var);
      mul_224 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_228_inst
    process(mul_224, conv65_219) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_224, conv65_219, tmp_var);
      mul66_229 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_272_inst
    process(conv84_260, conv82_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_260, conv82_256, tmp_var);
      mul85_273 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_277_inst
    process(mul85_273, conv87_264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_273, conv87_264, tmp_var);
      mul88_278 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_282_inst
    process(mul88_278, conv90_268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_278, conv90_268, tmp_var);
      mul91_283 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_863_inst
    process(conv255_855, conv253_851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_855, conv253_851, tmp_var);
      mul256_864 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_868_inst
    process(mul256_864, conv258_859) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_864, conv258_859, tmp_var);
      mul259_869 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_106_inst
    process(shl18_95, conv20_102) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_95, conv20_102, tmp_var);
      add21_107 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_131_inst
    process(shl27_120, conv29_127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_120, conv29_127, tmp_var);
      add30_132 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_156_inst
    process(shl36_145, conv38_152) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_145, conv38_152, tmp_var);
      add39_157 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_181_inst
    process(shl45_170, conv47_177) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_170, conv47_177, tmp_var);
      add48_182 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_206_inst
    process(shl54_195, conv56_202) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_195, conv56_202, tmp_var);
      add57_207 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_307_inst
    process(shl96_296, conv98_303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_296, conv98_303, tmp_var);
      add99_308 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_332_inst
    process(shl105_321, conv107_328) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_321, conv107_328, tmp_var);
      add108_333 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_357_inst
    process(shl114_346, conv116_353) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_346, conv116_353, tmp_var);
      add117_358 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_382_inst
    process(shl123_371, conv125_378) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_371, conv125_378, tmp_var);
      add126_383 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_407_inst
    process(shl132_396, conv134_403) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_396, conv134_403, tmp_var);
      add135_408 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_56_inst
    process(shl_45, conv3_52) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_45, conv3_52, tmp_var);
      add_57 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_81_inst
    process(shl9_70, conv11_77) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_70, conv11_77, tmp_var);
      add12_82 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_507_inst
    process(shl146_496, conv149_503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_496, conv149_503, tmp_var);
      add150_508 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_525_inst
    process(shl152_514, conv155_521) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_514, conv155_521, tmp_var);
      add156_526 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_543_inst
    process(shl158_532, conv161_539) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_532, conv161_539, tmp_var);
      add162_544 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_561_inst
    process(shl164_550, conv167_557) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_550, conv167_557, tmp_var);
      add168_562 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_579_inst
    process(shl170_568, conv173_575) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_568, conv173_575, tmp_var);
      add174_580 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_597_inst
    process(shl176_586, conv179_593) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_586, conv179_593, tmp_var);
      add180_598 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_615_inst
    process(shl182_604, conv185_611) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_604, conv185_611, tmp_var);
      add186_616 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_714_inst
    process(shl202_703, conv205_710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_703, conv205_710, tmp_var);
      add206_715 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_732_inst
    process(shl208_721, conv211_728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_721, conv211_728, tmp_var);
      add212_733 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_750_inst
    process(shl214_739, conv217_746) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_739, conv217_746, tmp_var);
      add218_751 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_768_inst
    process(shl220_757, conv223_764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_757, conv223_764, tmp_var);
      add224_769 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_786_inst
    process(shl226_775, conv229_782) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_775, conv229_782, tmp_var);
      add230_787 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_804_inst
    process(shl232_793, conv235_800) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_793, conv235_800, tmp_var);
      add236_805 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_822_inst
    process(shl238_811, conv241_818) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_811, conv241_818, tmp_var);
      add242_823 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_119_inst
    process(conv26_114) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_114, type_cast_118_wire_constant, tmp_var);
      shl27_120 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_144_inst
    process(conv35_139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_139, type_cast_143_wire_constant, tmp_var);
      shl36_145 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_169_inst
    process(conv44_164) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_164, type_cast_168_wire_constant, tmp_var);
      shl45_170 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_194_inst
    process(conv53_189) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_189, type_cast_193_wire_constant, tmp_var);
      shl54_195 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_295_inst
    process(conv95_290) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_290, type_cast_294_wire_constant, tmp_var);
      shl96_296 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_320_inst
    process(conv104_315) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_315, type_cast_319_wire_constant, tmp_var);
      shl105_321 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_345_inst
    process(conv113_340) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_340, type_cast_344_wire_constant, tmp_var);
      shl114_346 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_370_inst
    process(conv122_365) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_365, type_cast_369_wire_constant, tmp_var);
      shl123_371 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_395_inst
    process(conv131_390) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_390, type_cast_394_wire_constant, tmp_var);
      shl132_396 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_44_inst
    process(conv1_39) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_39, type_cast_43_wire_constant, tmp_var);
      shl_45 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_69_inst
    process(conv8_64) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_64, type_cast_68_wire_constant, tmp_var);
      shl9_70 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_94_inst
    process(conv17_89) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_89, type_cast_93_wire_constant, tmp_var);
      shl18_95 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_495_inst
    process(conv144_490) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_490, type_cast_494_wire_constant, tmp_var);
      shl146_496 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_513_inst
    process(add150_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_508, type_cast_512_wire_constant, tmp_var);
      shl152_514 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_531_inst
    process(add156_526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_526, type_cast_530_wire_constant, tmp_var);
      shl158_532 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_549_inst
    process(add162_544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_544, type_cast_548_wire_constant, tmp_var);
      shl164_550 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_567_inst
    process(add168_562) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_562, type_cast_566_wire_constant, tmp_var);
      shl170_568 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_585_inst
    process(add174_580) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_580, type_cast_584_wire_constant, tmp_var);
      shl176_586 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_603_inst
    process(add180_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_598, type_cast_602_wire_constant, tmp_var);
      shl182_604 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_702_inst
    process(conv200_697) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_697, type_cast_701_wire_constant, tmp_var);
      shl202_703 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_720_inst
    process(add206_715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_715, type_cast_719_wire_constant, tmp_var);
      shl208_721 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_738_inst
    process(add212_733) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_733, type_cast_737_wire_constant, tmp_var);
      shl214_739 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_756_inst
    process(add218_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_751, type_cast_755_wire_constant, tmp_var);
      shl220_757 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_774_inst
    process(add224_769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_769, type_cast_773_wire_constant, tmp_var);
      shl226_775 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_792_inst
    process(add230_787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_787, type_cast_791_wire_constant, tmp_var);
      shl232_793 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_810_inst
    process(add236_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_805, type_cast_809_wire_constant, tmp_var);
      shl238_811 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1205_inst
    process(conv355_1201, conv276_968) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1201, conv276_968, tmp_var);
      sub_1206 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1323_inst
    process(tmp520_1318) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp520_1318, type_cast_1322_wire_constant, tmp_var);
      tmp521_1324 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_413_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_229, type_cast_412_wire_constant, tmp_var);
      cmp513_415 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_429_inst
    process(mul91_283) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_283, type_cast_428_wire_constant, tmp_var);
      cmp194509_430 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_442_inst
    process(shr_235) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_235, type_cast_441_wire_constant, tmp_var);
      tmp563_443 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_649_inst
    process(tmp548_644) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp548_644, type_cast_648_wire_constant, tmp_var);
      tmp549_650 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_874_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_869, type_cast_873_wire_constant, tmp_var);
      cmp264505_875 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_893_inst
    process(tmp532_888) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp532_888, type_cast_892_wire_constant, tmp_var);
      tmp533_894 <= tmp_var; --
    end process;
    -- shared split operator group (107) : array_obj_ref_1362_index_offset 
    ApIntAdd_group_107: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1361_scaled;
      array_obj_ref_1362_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1362_index_offset_req_0;
      array_obj_ref_1362_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1362_index_offset_req_1;
      array_obj_ref_1362_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_107_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_107_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_107",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : array_obj_ref_481_index_offset 
    ApIntAdd_group_108: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar555_480_scaled;
      array_obj_ref_481_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_481_index_offset_req_0;
      array_obj_ref_481_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_481_index_offset_req_1;
      array_obj_ref_481_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_108_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_108_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_108",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : array_obj_ref_688_index_offset 
    ApIntAdd_group_109: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar539_687_scaled;
      array_obj_ref_688_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_688_index_offset_req_0;
      array_obj_ref_688_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_688_index_offset_req_1;
      array_obj_ref_688_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_109_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_109_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : array_obj_ref_932_index_offset 
    ApIntAdd_group_110: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar525_931_scaled;
      array_obj_ref_932_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_932_index_offset_req_0;
      array_obj_ref_932_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_932_index_offset_req_1;
      array_obj_ref_932_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_110_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_110_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- unary operator type_cast_1199_inst
    process(call354_1196) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1196, tmp_var);
      type_cast_1199_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_966_inst
    process(call275_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_962, tmp_var);
      type_cast_966_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1367_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1367_load_0_req_0;
      ptr_deref_1367_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1367_load_0_req_1;
      ptr_deref_1367_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1367_word_address_0;
      ptr_deref_1367_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_618_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_618_store_0_req_0;
      ptr_deref_618_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_618_store_0_req_1;
      ptr_deref_618_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_618_word_address_0;
      data_in <= ptr_deref_618_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_825_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_825_store_0_req_0;
      ptr_deref_825_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_825_store_0_req_1;
      ptr_deref_825_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_825_word_address_0;
      data_in <= ptr_deref_825_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_936_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_936_store_0_req_0;
      ptr_deref_936_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_936_store_0_req_1;
      ptr_deref_936_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_936_word_address_0;
      data_in <= ptr_deref_936_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1183_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1183_inst_req_0;
      RPIPE_Block0_done_1183_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1183_inst_req_1;
      RPIPE_Block0_done_1183_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1184 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1186_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1186_inst_req_0;
      RPIPE_Block1_done_1186_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1186_inst_req_1;
      RPIPE_Block1_done_1186_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1187 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1189_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1189_inst_req_0;
      RPIPE_Block2_done_1189_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1189_inst_req_1;
      RPIPE_Block2_done_1189_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1190 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1192_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1192_inst_req_0;
      RPIPE_Block3_done_1192_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1192_inst_req_1;
      RPIPE_Block3_done_1192_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1193 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_759_inst RPIPE_ConvTranspose_input_pipe_59_inst RPIPE_ConvTranspose_input_pipe_84_inst RPIPE_ConvTranspose_input_pipe_741_inst RPIPE_ConvTranspose_input_pipe_47_inst RPIPE_ConvTranspose_input_pipe_97_inst RPIPE_ConvTranspose_input_pipe_147_inst RPIPE_ConvTranspose_input_pipe_122_inst RPIPE_ConvTranspose_input_pipe_777_inst RPIPE_ConvTranspose_input_pipe_159_inst RPIPE_ConvTranspose_input_pipe_795_inst RPIPE_ConvTranspose_input_pipe_134_inst RPIPE_ConvTranspose_input_pipe_692_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_813_inst RPIPE_ConvTranspose_input_pipe_109_inst RPIPE_ConvTranspose_input_pipe_705_inst RPIPE_ConvTranspose_input_pipe_172_inst RPIPE_ConvTranspose_input_pipe_72_inst RPIPE_ConvTranspose_input_pipe_723_inst RPIPE_ConvTranspose_input_pipe_184_inst RPIPE_ConvTranspose_input_pipe_197_inst RPIPE_ConvTranspose_input_pipe_285_inst RPIPE_ConvTranspose_input_pipe_298_inst RPIPE_ConvTranspose_input_pipe_310_inst RPIPE_ConvTranspose_input_pipe_323_inst RPIPE_ConvTranspose_input_pipe_335_inst RPIPE_ConvTranspose_input_pipe_348_inst RPIPE_ConvTranspose_input_pipe_360_inst RPIPE_ConvTranspose_input_pipe_373_inst RPIPE_ConvTranspose_input_pipe_385_inst RPIPE_ConvTranspose_input_pipe_398_inst RPIPE_ConvTranspose_input_pipe_485_inst RPIPE_ConvTranspose_input_pipe_498_inst RPIPE_ConvTranspose_input_pipe_516_inst RPIPE_ConvTranspose_input_pipe_534_inst RPIPE_ConvTranspose_input_pipe_552_inst RPIPE_ConvTranspose_input_pipe_570_inst RPIPE_ConvTranspose_input_pipe_588_inst RPIPE_ConvTranspose_input_pipe_606_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_692_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_813_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_285_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_298_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_310_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_323_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_335_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_348_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_360_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_373_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_385_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_398_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_485_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_498_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_516_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_552_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_570_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_588_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_606_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_692_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_813_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_285_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_298_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_310_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_323_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_335_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_348_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_360_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_373_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_385_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_398_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_485_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_498_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_516_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_552_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_570_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_588_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_606_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_692_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_813_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_285_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_298_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_310_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_323_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_335_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_348_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_360_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_373_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_385_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_398_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_485_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_498_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_516_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_552_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_570_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_588_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_606_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_692_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_813_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_285_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_298_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_310_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_323_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_335_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_348_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_360_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_373_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_385_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_398_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_485_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_498_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_516_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_552_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_570_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_588_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_606_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call221_760 <= data_out(319 downto 312);
      call5_60 <= data_out(311 downto 304);
      call14_85 <= data_out(303 downto 296);
      call215_742 <= data_out(295 downto 288);
      call2_48 <= data_out(287 downto 280);
      call19_98 <= data_out(279 downto 272);
      call37_148 <= data_out(271 downto 264);
      call28_123 <= data_out(263 downto 256);
      call227_778 <= data_out(255 downto 248);
      call41_160 <= data_out(247 downto 240);
      call233_796 <= data_out(239 downto 232);
      call32_135 <= data_out(231 downto 224);
      call199_693 <= data_out(223 downto 216);
      call_35 <= data_out(215 downto 208);
      call239_814 <= data_out(207 downto 200);
      call23_110 <= data_out(199 downto 192);
      call203_706 <= data_out(191 downto 184);
      call46_173 <= data_out(183 downto 176);
      call10_73 <= data_out(175 downto 168);
      call209_724 <= data_out(167 downto 160);
      call50_185 <= data_out(159 downto 152);
      call55_198 <= data_out(151 downto 144);
      call92_286 <= data_out(143 downto 136);
      call97_299 <= data_out(135 downto 128);
      call101_311 <= data_out(127 downto 120);
      call106_324 <= data_out(119 downto 112);
      call110_336 <= data_out(111 downto 104);
      call115_349 <= data_out(103 downto 96);
      call119_361 <= data_out(95 downto 88);
      call124_374 <= data_out(87 downto 80);
      call128_386 <= data_out(79 downto 72);
      call133_399 <= data_out(71 downto 64);
      call143_486 <= data_out(63 downto 56);
      call147_499 <= data_out(55 downto 48);
      call153_517 <= data_out(47 downto 40);
      call159_535 <= data_out(39 downto 32);
      call165_553 <= data_out(31 downto 24);
      call171_571 <= data_out(23 downto 16);
      call177_589 <= data_out(15 downto 8);
      call183_607 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_1008_inst WPIPE_Block0_start_997_inst WPIPE_Block0_start_1011_inst WPIPE_Block0_start_970_inst WPIPE_Block0_start_973_inst WPIPE_Block0_start_976_inst WPIPE_Block0_start_1001_inst WPIPE_Block0_start_979_inst WPIPE_Block0_start_982_inst WPIPE_Block0_start_1005_inst WPIPE_Block0_start_985_inst WPIPE_Block0_start_988_inst WPIPE_Block0_start_991_inst WPIPE_Block0_start_994_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_1008_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_997_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_1011_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_970_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_973_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_976_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_1001_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_979_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_982_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_1005_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_985_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_988_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_991_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_994_inst_req_0;
      WPIPE_Block0_start_1008_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_997_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_1011_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_970_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_973_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_976_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_1001_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_979_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_982_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_1005_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_985_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_988_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_991_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_994_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_1008_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_997_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_1011_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_970_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_973_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_976_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_1001_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_979_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_982_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_1005_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_985_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_988_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_991_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_994_inst_req_1;
      WPIPE_Block0_start_1008_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_997_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_1011_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_970_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_973_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_976_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_1001_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_979_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_982_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_1005_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_985_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_988_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_991_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_994_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add126_383 & type_cast_999_wire_constant & add135_408 & add_57 & add12_82 & add21_107 & type_cast_1003_wire_constant & add30_132 & add39_157 & add117_358 & add48_182 & add57_207 & add99_308 & add108_333;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1051_inst WPIPE_Block1_start_1067_inst WPIPE_Block1_start_1064_inst WPIPE_Block1_start_1061_inst WPIPE_Block1_start_1058_inst WPIPE_Block1_start_1014_inst WPIPE_Block1_start_1017_inst WPIPE_Block1_start_1020_inst WPIPE_Block1_start_1023_inst WPIPE_Block1_start_1026_inst WPIPE_Block1_start_1029_inst WPIPE_Block1_start_1032_inst WPIPE_Block1_start_1035_inst WPIPE_Block1_start_1038_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1051_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1067_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1064_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1061_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1058_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1014_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1017_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1020_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1023_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1026_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1029_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1032_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1035_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1038_inst_req_0;
      WPIPE_Block1_start_1051_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1067_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1064_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1061_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1058_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1014_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1017_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1020_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1023_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1026_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1029_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1032_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1035_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1038_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1051_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1067_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1064_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1061_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1058_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1014_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1017_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1020_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1023_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1026_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1029_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1032_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1035_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1038_inst_req_1;
      WPIPE_Block1_start_1051_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1067_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1064_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1061_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1058_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1014_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1017_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1020_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1023_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1026_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1029_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1032_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1035_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1038_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= conv305_1050 & add135_408 & add126_383 & add117_358 & conv307_1057 & add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_308 & add108_333;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1114_inst WPIPE_Block2_start_1123_inst WPIPE_Block2_start_1120_inst WPIPE_Block2_start_1070_inst WPIPE_Block2_start_1073_inst WPIPE_Block2_start_1076_inst WPIPE_Block2_start_1117_inst WPIPE_Block2_start_1079_inst WPIPE_Block2_start_1082_inst WPIPE_Block2_start_1085_inst WPIPE_Block2_start_1088_inst WPIPE_Block2_start_1091_inst WPIPE_Block2_start_1094_inst WPIPE_Block2_start_1107_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1114_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1123_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1120_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1070_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1073_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1076_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1117_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1079_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1082_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1085_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1088_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1091_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1094_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1107_inst_req_0;
      WPIPE_Block2_start_1114_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1123_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1120_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1070_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1073_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1076_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1117_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1079_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1082_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1085_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1088_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1091_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1094_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1107_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1114_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1123_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1120_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1070_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1073_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1076_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1117_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1079_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1082_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1085_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1088_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1091_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1094_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1107_inst_req_1;
      WPIPE_Block2_start_1114_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1123_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1120_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1070_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1073_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1076_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1117_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1079_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1082_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1085_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1088_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1091_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1094_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1107_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= conv324_1113 & add135_408 & add126_383 & add_57 & add12_82 & add21_107 & add117_358 & add30_132 & add39_157 & add48_182 & add57_207 & add99_308 & add108_333 & conv322_1106;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1126_inst WPIPE_Block3_start_1176_inst WPIPE_Block3_start_1129_inst WPIPE_Block3_start_1132_inst WPIPE_Block3_start_1135_inst WPIPE_Block3_start_1141_inst WPIPE_Block3_start_1179_inst WPIPE_Block3_start_1144_inst WPIPE_Block3_start_1170_inst WPIPE_Block3_start_1150_inst WPIPE_Block3_start_1163_inst WPIPE_Block3_start_1173_inst WPIPE_Block3_start_1138_inst WPIPE_Block3_start_1147_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1126_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1176_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1129_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1132_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1135_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1141_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1179_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1144_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1170_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1150_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1163_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1173_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1138_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1147_inst_req_0;
      WPIPE_Block3_start_1126_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1176_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1129_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1132_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1135_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1141_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1179_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1144_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1170_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1150_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1163_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1173_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1138_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1147_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1126_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1176_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1129_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1132_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1135_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1141_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1179_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1144_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1170_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1150_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1163_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1173_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1138_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1147_inst_req_1;
      WPIPE_Block3_start_1126_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1176_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1129_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1132_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1135_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1141_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1179_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1144_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1170_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1150_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1163_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1173_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1138_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1147_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add_57 & add126_383 & add12_82 & add21_107 & add30_132 & add48_182 & add135_408 & add57_207 & conv341_1169 & add108_333 & conv339_1162 & add117_358 & add39_157 & add99_308;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1284_inst WPIPE_ConvTranspose_output_pipe_1299_inst WPIPE_ConvTranspose_output_pipe_1287_inst WPIPE_ConvTranspose_output_pipe_1281_inst WPIPE_ConvTranspose_output_pipe_1290_inst WPIPE_ConvTranspose_output_pipe_1302_inst WPIPE_ConvTranspose_output_pipe_1296_inst WPIPE_ConvTranspose_output_pipe_1293_inst WPIPE_ConvTranspose_output_pipe_1443_inst WPIPE_ConvTranspose_output_pipe_1446_inst WPIPE_ConvTranspose_output_pipe_1449_inst WPIPE_ConvTranspose_output_pipe_1452_inst WPIPE_ConvTranspose_output_pipe_1455_inst WPIPE_ConvTranspose_output_pipe_1458_inst WPIPE_ConvTranspose_output_pipe_1461_inst WPIPE_ConvTranspose_output_pipe_1464_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1284_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1299_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1281_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1302_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1296_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1293_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1443_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1446_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1449_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1452_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1455_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1458_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1461_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1464_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1443_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1446_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1284_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1299_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1281_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1302_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1296_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1293_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1443_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1446_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1449_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1452_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1455_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1458_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1461_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1464_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1443_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1446_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv397_1270 & conv367_1220 & conv391_1260 & conv403_1280 & conv385_1250 & conv361_1210 & conv373_1230 & conv379_1240 & conv479_1442 & conv473_1432 & conv467_1422 & conv461_1412 & conv455_1402 & conv449_1392 & conv443_1382 & conv437_1372;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1196_call call_stmt_962_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1196_call_req_0;
      reqL_unguarded(0) <= call_stmt_962_call_req_0;
      call_stmt_1196_call_ack_0 <= ackL_unguarded(1);
      call_stmt_962_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1196_call_req_1;
      reqR_unguarded(0) <= call_stmt_962_call_req_1;
      call_stmt_1196_call_ack_1 <= ackR_unguarded(1);
      call_stmt_962_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call354_1196 <= data_out(127 downto 64);
      call275_962 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3763_start: Boolean;
  signal convTransposeA_CP_3763_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1826_inst_req_1 : boolean;
  signal type_cast_1816_inst_ack_1 : boolean;
  signal type_cast_1621_inst_req_1 : boolean;
  signal type_cast_1621_inst_ack_1 : boolean;
  signal type_cast_1822_inst_req_0 : boolean;
  signal phi_stmt_1817_req_1 : boolean;
  signal type_cast_1822_inst_req_1 : boolean;
  signal type_cast_1614_inst_req_0 : boolean;
  signal type_cast_1607_inst_req_0 : boolean;
  signal phi_stmt_1810_ack_0 : boolean;
  signal type_cast_1822_inst_ack_0 : boolean;
  signal type_cast_1816_inst_req_1 : boolean;
  signal phi_stmt_1615_req_0 : boolean;
  signal phi_stmt_1810_req_1 : boolean;
  signal phi_stmt_1615_req_1 : boolean;
  signal type_cast_1607_inst_req_1 : boolean;
  signal type_cast_1614_inst_req_1 : boolean;
  signal type_cast_1607_inst_ack_0 : boolean;
  signal type_cast_1614_inst_ack_1 : boolean;
  signal phi_stmt_1601_req_1 : boolean;
  signal type_cast_1607_inst_ack_1 : boolean;
  signal phi_stmt_1823_req_0 : boolean;
  signal type_cast_1614_inst_ack_0 : boolean;
  signal phi_stmt_1608_req_1 : boolean;
  signal type_cast_1822_inst_ack_1 : boolean;
  signal type_cast_1621_inst_ack_0 : boolean;
  signal type_cast_1826_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1497_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1503_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1506_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1506_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1512_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1506_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1506_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1500_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1500_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1509_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1509_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1512_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1503_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1497_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1497_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1503_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1494_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1494_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1500_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1494_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1503_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1512_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1512_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1500_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1497_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1494_inst_ack_1 : boolean;
  signal phi_stmt_1622_req_0 : boolean;
  signal phi_stmt_1817_ack_0 : boolean;
  signal type_cast_1828_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1515_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1515_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1515_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1515_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1518_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1518_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1518_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1518_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1521_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1521_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1521_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1521_inst_ack_1 : boolean;
  signal type_cast_1525_inst_req_0 : boolean;
  signal type_cast_1525_inst_ack_0 : boolean;
  signal type_cast_1525_inst_req_1 : boolean;
  signal type_cast_1525_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1534_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1534_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1534_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1534_inst_ack_1 : boolean;
  signal type_cast_1538_inst_req_0 : boolean;
  signal type_cast_1538_inst_ack_0 : boolean;
  signal type_cast_1538_inst_req_1 : boolean;
  signal type_cast_1538_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1546_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1546_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1546_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1546_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1549_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1549_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1549_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1549_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1552_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1552_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1552_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1552_inst_ack_1 : boolean;
  signal phi_stmt_1823_ack_0 : boolean;
  signal type_cast_1579_inst_req_0 : boolean;
  signal type_cast_1579_inst_ack_0 : boolean;
  signal type_cast_1579_inst_req_1 : boolean;
  signal type_cast_1579_inst_ack_1 : boolean;
  signal type_cast_1583_inst_req_0 : boolean;
  signal type_cast_1583_inst_ack_0 : boolean;
  signal type_cast_1583_inst_req_1 : boolean;
  signal type_cast_1583_inst_ack_1 : boolean;
  signal type_cast_1587_inst_req_0 : boolean;
  signal type_cast_1587_inst_ack_0 : boolean;
  signal type_cast_1587_inst_req_1 : boolean;
  signal type_cast_1587_inst_ack_1 : boolean;
  signal type_cast_1591_inst_req_0 : boolean;
  signal type_cast_1591_inst_ack_0 : boolean;
  signal type_cast_1591_inst_req_1 : boolean;
  signal type_cast_1591_inst_ack_1 : boolean;
  signal type_cast_1663_inst_req_0 : boolean;
  signal type_cast_1663_inst_ack_0 : boolean;
  signal type_cast_1663_inst_req_1 : boolean;
  signal type_cast_1663_inst_ack_1 : boolean;
  signal type_cast_1667_inst_req_0 : boolean;
  signal type_cast_1667_inst_ack_0 : boolean;
  signal type_cast_1667_inst_req_1 : boolean;
  signal type_cast_1667_inst_ack_1 : boolean;
  signal type_cast_1671_inst_req_0 : boolean;
  signal type_cast_1671_inst_ack_0 : boolean;
  signal type_cast_1671_inst_req_1 : boolean;
  signal type_cast_1671_inst_ack_1 : boolean;
  signal type_cast_1701_inst_req_0 : boolean;
  signal type_cast_1701_inst_ack_0 : boolean;
  signal type_cast_1701_inst_req_1 : boolean;
  signal type_cast_1701_inst_ack_1 : boolean;
  signal type_cast_1621_inst_req_0 : boolean;
  signal phi_stmt_1608_req_0 : boolean;
  signal type_cast_1826_inst_ack_0 : boolean;
  signal type_cast_1826_inst_req_0 : boolean;
  signal array_obj_ref_1707_index_offset_req_0 : boolean;
  signal phi_stmt_1810_req_0 : boolean;
  signal array_obj_ref_1707_index_offset_ack_0 : boolean;
  signal array_obj_ref_1707_index_offset_req_1 : boolean;
  signal array_obj_ref_1707_index_offset_ack_1 : boolean;
  signal addr_of_1708_final_reg_req_0 : boolean;
  signal addr_of_1708_final_reg_ack_0 : boolean;
  signal addr_of_1708_final_reg_req_1 : boolean;
  signal addr_of_1708_final_reg_ack_1 : boolean;
  signal phi_stmt_1823_req_1 : boolean;
  signal type_cast_1828_inst_ack_1 : boolean;
  signal type_cast_1828_inst_req_1 : boolean;
  signal phi_stmt_1817_req_0 : boolean;
  signal ptr_deref_1712_load_0_req_0 : boolean;
  signal ptr_deref_1712_load_0_ack_0 : boolean;
  signal ptr_deref_1712_load_0_req_1 : boolean;
  signal ptr_deref_1712_load_0_ack_1 : boolean;
  signal type_cast_1816_inst_ack_0 : boolean;
  signal phi_stmt_1622_ack_0 : boolean;
  signal phi_stmt_1615_ack_0 : boolean;
  signal phi_stmt_1608_ack_0 : boolean;
  signal phi_stmt_1601_ack_0 : boolean;
  signal phi_stmt_1622_req_1 : boolean;
  signal type_cast_1628_inst_ack_1 : boolean;
  signal type_cast_1628_inst_req_1 : boolean;
  signal type_cast_1628_inst_ack_0 : boolean;
  signal array_obj_ref_1730_index_offset_req_0 : boolean;
  signal type_cast_1820_inst_ack_1 : boolean;
  signal array_obj_ref_1730_index_offset_ack_0 : boolean;
  signal array_obj_ref_1730_index_offset_req_1 : boolean;
  signal type_cast_1820_inst_req_1 : boolean;
  signal array_obj_ref_1730_index_offset_ack_1 : boolean;
  signal type_cast_1816_inst_req_0 : boolean;
  signal type_cast_1628_inst_req_0 : boolean;
  signal addr_of_1731_final_reg_req_0 : boolean;
  signal type_cast_1820_inst_ack_0 : boolean;
  signal addr_of_1731_final_reg_ack_0 : boolean;
  signal addr_of_1731_final_reg_req_1 : boolean;
  signal type_cast_1820_inst_req_0 : boolean;
  signal addr_of_1731_final_reg_ack_1 : boolean;
  signal type_cast_1828_inst_ack_0 : boolean;
  signal ptr_deref_1734_store_0_req_0 : boolean;
  signal ptr_deref_1734_store_0_ack_0 : boolean;
  signal ptr_deref_1734_store_0_req_1 : boolean;
  signal ptr_deref_1734_store_0_ack_1 : boolean;
  signal type_cast_1739_inst_req_0 : boolean;
  signal type_cast_1739_inst_ack_0 : boolean;
  signal type_cast_1739_inst_req_1 : boolean;
  signal type_cast_1739_inst_ack_1 : boolean;
  signal if_stmt_1752_branch_req_0 : boolean;
  signal if_stmt_1752_branch_ack_1 : boolean;
  signal if_stmt_1752_branch_ack_0 : boolean;
  signal type_cast_1780_inst_req_0 : boolean;
  signal type_cast_1780_inst_ack_0 : boolean;
  signal type_cast_1780_inst_req_1 : boolean;
  signal type_cast_1780_inst_ack_1 : boolean;
  signal type_cast_1796_inst_req_0 : boolean;
  signal type_cast_1796_inst_ack_0 : boolean;
  signal type_cast_1796_inst_req_1 : boolean;
  signal type_cast_1796_inst_ack_1 : boolean;
  signal if_stmt_1803_branch_req_0 : boolean;
  signal if_stmt_1803_branch_ack_1 : boolean;
  signal if_stmt_1803_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1839_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1839_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1839_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1839_inst_ack_1 : boolean;
  signal phi_stmt_1601_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3763_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3763: Block -- control-path 
    signal convTransposeA_CP_3763_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3763_elements(0) <= convTransposeA_CP_3763_start;
    convTransposeA_CP_3763_symbol <= convTransposeA_CP_3763_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1492/branch_block_stmt_1492__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553__entry__
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/$entry
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1492/$entry
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_Update/cr
      -- 
    rr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => RPIPE_Block0_start_1494_inst_req_0); -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => type_cast_1525_inst_req_1); -- 
    cr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => type_cast_1538_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/merge_stmt_1809__exit__
      -- CP-element group 1: 	 branch_block_stmt_1492/assign_stmt_1835__entry__
      -- CP-element group 1: 	 branch_block_stmt_1492/assign_stmt_1835__exit__
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/assign_stmt_1835/$entry
      -- CP-element group 1: 	 branch_block_stmt_1492/assign_stmt_1835/$exit
      -- 
    cr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1621_inst_req_1); -- 
    rr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1614_inst_req_0); -- 
    rr_4497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1607_inst_req_0); -- 
    cr_4502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1607_inst_req_1); -- 
    cr_4525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1614_inst_req_1); -- 
    rr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1621_inst_req_0); -- 
    cr_4571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1628_inst_req_1); -- 
    rr_4566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => type_cast_1628_inst_req_0); -- 
    convTransposeA_CP_3763_elements(1) <= convTransposeA_CP_3763_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_Update/cr
      -- 
    ra_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1494_inst_ack_0, ack => convTransposeA_CP_3763_elements(2)); -- 
    cr_3816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(2), ack => RPIPE_Block0_start_1494_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1494_Update/ca
      -- 
    ca_3817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1494_inst_ack_1, ack => convTransposeA_CP_3763_elements(3)); -- 
    rr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(3), ack => RPIPE_Block0_start_1497_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_Update/$entry
      -- 
    ra_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1497_inst_ack_0, ack => convTransposeA_CP_3763_elements(4)); -- 
    cr_3830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(4), ack => RPIPE_Block0_start_1497_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1497_Update/ca
      -- 
    ca_3831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1497_inst_ack_1, ack => convTransposeA_CP_3763_elements(5)); -- 
    rr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(5), ack => RPIPE_Block0_start_1500_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_Sample/ra
      -- 
    ra_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1500_inst_ack_0, ack => convTransposeA_CP_3763_elements(6)); -- 
    cr_3844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(6), ack => RPIPE_Block0_start_1500_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1500_update_completed_
      -- 
    ca_3845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1500_inst_ack_1, ack => convTransposeA_CP_3763_elements(7)); -- 
    rr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(7), ack => RPIPE_Block0_start_1503_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_Update/cr
      -- 
    ra_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1503_inst_ack_0, ack => convTransposeA_CP_3763_elements(8)); -- 
    cr_3858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(8), ack => RPIPE_Block0_start_1503_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1503_Update/$exit
      -- 
    ca_3859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1503_inst_ack_1, ack => convTransposeA_CP_3763_elements(9)); -- 
    rr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(9), ack => RPIPE_Block0_start_1506_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_Update/$entry
      -- 
    ra_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1506_inst_ack_0, ack => convTransposeA_CP_3763_elements(10)); -- 
    cr_3872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(10), ack => RPIPE_Block0_start_1506_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1506_update_completed_
      -- 
    ca_3873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1506_inst_ack_1, ack => convTransposeA_CP_3763_elements(11)); -- 
    rr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(11), ack => RPIPE_Block0_start_1509_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_sample_completed_
      -- 
    ra_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1509_inst_ack_0, ack => convTransposeA_CP_3763_elements(12)); -- 
    cr_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(12), ack => RPIPE_Block0_start_1509_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1509_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_Sample/rr
      -- 
    ca_3887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1509_inst_ack_1, ack => convTransposeA_CP_3763_elements(13)); -- 
    rr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(13), ack => RPIPE_Block0_start_1512_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_Sample/ra
      -- 
    ra_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1512_inst_ack_0, ack => convTransposeA_CP_3763_elements(14)); -- 
    cr_3900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(14), ack => RPIPE_Block0_start_1512_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1512_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_Sample/rr
      -- 
    ca_3901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1512_inst_ack_1, ack => convTransposeA_CP_3763_elements(15)); -- 
    rr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(15), ack => RPIPE_Block0_start_1515_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_Update/cr
      -- 
    ra_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1515_inst_ack_0, ack => convTransposeA_CP_3763_elements(16)); -- 
    cr_3914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(16), ack => RPIPE_Block0_start_1515_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1515_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_Sample/rr
      -- 
    ca_3915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1515_inst_ack_1, ack => convTransposeA_CP_3763_elements(17)); -- 
    rr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(17), ack => RPIPE_Block0_start_1518_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_Update/cr
      -- 
    ra_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1518_inst_ack_0, ack => convTransposeA_CP_3763_elements(18)); -- 
    cr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(18), ack => RPIPE_Block0_start_1518_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1518_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_Sample/rr
      -- 
    ca_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1518_inst_ack_1, ack => convTransposeA_CP_3763_elements(19)); -- 
    rr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(19), ack => RPIPE_Block0_start_1521_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_Update/cr
      -- 
    ra_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1521_inst_ack_0, ack => convTransposeA_CP_3763_elements(20)); -- 
    cr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(20), ack => RPIPE_Block0_start_1521_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1521_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_Sample/rr
      -- 
    ca_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1521_inst_ack_1, ack => convTransposeA_CP_3763_elements(21)); -- 
    rr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(21), ack => type_cast_1525_inst_req_0); -- 
    rr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(21), ack => RPIPE_Block0_start_1534_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_Sample/ra
      -- 
    ra_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1525_inst_ack_0, ack => convTransposeA_CP_3763_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1525_Update/ca
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1525_inst_ack_1, ack => convTransposeA_CP_3763_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_Update/cr
      -- 
    ra_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1534_inst_ack_0, ack => convTransposeA_CP_3763_elements(24)); -- 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(24), ack => RPIPE_Block0_start_1534_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1534_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_Sample/rr
      -- 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1534_inst_ack_1, ack => convTransposeA_CP_3763_elements(25)); -- 
    rr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(25), ack => type_cast_1538_inst_req_0); -- 
    rr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(25), ack => RPIPE_Block0_start_1546_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_Sample/ra
      -- 
    ra_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_0, ack => convTransposeA_CP_3763_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/type_cast_1538_Update/ca
      -- 
    ca_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_1, ack => convTransposeA_CP_3763_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_Update/cr
      -- 
    ra_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1546_inst_ack_0, ack => convTransposeA_CP_3763_elements(28)); -- 
    cr_3998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(28), ack => RPIPE_Block0_start_1546_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1546_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_Sample/rr
      -- 
    ca_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1546_inst_ack_1, ack => convTransposeA_CP_3763_elements(29)); -- 
    rr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(29), ack => RPIPE_Block0_start_1549_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_Update/cr
      -- 
    ra_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1549_inst_ack_0, ack => convTransposeA_CP_3763_elements(30)); -- 
    cr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(30), ack => RPIPE_Block0_start_1549_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1549_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_Sample/rr
      -- 
    ca_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1549_inst_ack_1, ack => convTransposeA_CP_3763_elements(31)); -- 
    rr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(31), ack => RPIPE_Block0_start_1552_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_Update/cr
      -- 
    ra_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1552_inst_ack_0, ack => convTransposeA_CP_3763_elements(32)); -- 
    cr_4026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(32), ack => RPIPE_Block0_start_1552_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/RPIPE_Block0_start_1552_Update/ca
      -- 
    ca_4027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1552_inst_ack_1, ack => convTransposeA_CP_3763_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553__exit__
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598__entry__
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1495_to_assign_stmt_1553/$exit
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_Update/cr
      -- 
    rr_4038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1579_inst_req_0); -- 
    cr_4043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1579_inst_req_1); -- 
    rr_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1583_inst_req_0); -- 
    cr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1583_inst_req_1); -- 
    rr_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1587_inst_req_0); -- 
    cr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1587_inst_req_1); -- 
    rr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1591_inst_req_0); -- 
    cr_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1591_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(23) & convTransposeA_CP_3763_elements(27) & convTransposeA_CP_3763_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_Sample/ra
      -- 
    ra_4039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1579_inst_ack_0, ack => convTransposeA_CP_3763_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1579_Update/ca
      -- 
    ca_4044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1579_inst_ack_1, ack => convTransposeA_CP_3763_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_Sample/ra
      -- 
    ra_4053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1583_inst_ack_0, ack => convTransposeA_CP_3763_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1583_Update/ca
      -- 
    ca_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1583_inst_ack_1, ack => convTransposeA_CP_3763_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_Sample/ra
      -- 
    ra_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_0, ack => convTransposeA_CP_3763_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1587_Update/ca
      -- 
    ca_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_1, ack => convTransposeA_CP_3763_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_Sample/ra
      -- 
    ra_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1591_inst_ack_0, ack => convTransposeA_CP_3763_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/type_cast_1591_Update/ca
      -- 
    ca_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1591_inst_ack_1, ack => convTransposeA_CP_3763_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1622/$entry
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598__exit__
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1492/assign_stmt_1560_to_assign_stmt_1598/$exit
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1615/$entry
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1601/$entry
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1608/$entry
      -- CP-element group 43: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(36) & convTransposeA_CP_3763_elements(38) & convTransposeA_CP_3763_elements(40) & convTransposeA_CP_3763_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_Sample/ra
      -- 
    ra_4098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_0, ack => convTransposeA_CP_3763_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_Update/ca
      -- 
    ca_4103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_1, ack => convTransposeA_CP_3763_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_Sample/ra
      -- 
    ra_4112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_0, ack => convTransposeA_CP_3763_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_Update/ca
      -- 
    ca_4117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_1, ack => convTransposeA_CP_3763_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_Sample/ra
      -- 
    ra_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1671_inst_ack_0, ack => convTransposeA_CP_3763_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_Update/ca
      -- 
    ca_4131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1671_inst_ack_1, ack => convTransposeA_CP_3763_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_Sample/ra
      -- 
    ra_4140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_0, ack => convTransposeA_CP_3763_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_Sample/req
      -- 
    ca_4145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_1, ack => convTransposeA_CP_3763_elements(51)); -- 
    req_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(51), ack => array_obj_ref_1707_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_Sample/ack
      -- 
    ack_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1707_index_offset_ack_0, ack => convTransposeA_CP_3763_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_request/req
      -- 
    ack_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1707_index_offset_ack_1, ack => convTransposeA_CP_3763_elements(53)); -- 
    req_4185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(53), ack => addr_of_1708_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_request/ack
      -- 
    ack_4186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1708_final_reg_ack_0, ack => convTransposeA_CP_3763_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Sample/word_access_start/word_0/rr
      -- 
    ack_4191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1708_final_reg_ack_1, ack => convTransposeA_CP_3763_elements(55)); -- 
    rr_4224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(55), ack => ptr_deref_1712_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Sample/word_access_start/word_0/ra
      -- 
    ra_4225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1712_load_0_ack_0, ack => convTransposeA_CP_3763_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/ptr_deref_1712_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/ptr_deref_1712_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/ptr_deref_1712_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/ptr_deref_1712_Merge/merge_ack
      -- 
    ca_4236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1712_load_0_ack_1, ack => convTransposeA_CP_3763_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_Sample/req
      -- 
    req_4266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(58), ack => array_obj_ref_1730_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(45) & convTransposeA_CP_3763_elements(47) & convTransposeA_CP_3763_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_Sample/ack
      -- 
    ack_4267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1730_index_offset_ack_0, ack => convTransposeA_CP_3763_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_request/req
      -- 
    ack_4272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1730_index_offset_ack_1, ack => convTransposeA_CP_3763_elements(60)); -- 
    req_4281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(60), ack => addr_of_1731_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_request/ack
      -- 
    ack_4282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1731_final_reg_ack_0, ack => convTransposeA_CP_3763_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_word_addrgen/root_register_ack
      -- 
    ack_4287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1731_final_reg_ack_1, ack => convTransposeA_CP_3763_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/ptr_deref_1734_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/ptr_deref_1734_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/ptr_deref_1734_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/ptr_deref_1734_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/word_access_start/word_0/rr
      -- 
    rr_4325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(63), ack => ptr_deref_1734_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(57) & convTransposeA_CP_3763_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Sample/word_access_start/word_0/ra
      -- 
    ra_4326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1734_store_0_ack_0, ack => convTransposeA_CP_3763_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Update/word_access_complete/word_0/ca
      -- 
    ca_4337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1734_store_0_ack_1, ack => convTransposeA_CP_3763_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_Sample/ra
      -- 
    ra_4346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1739_inst_ack_0, ack => convTransposeA_CP_3763_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_Update/ca
      -- 
    ca_4351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1739_inst_ack_1, ack => convTransposeA_CP_3763_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751__exit__
      -- CP-element group 68: 	 branch_block_stmt_1492/if_stmt_1752__entry__
      -- CP-element group 68: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/$exit
      -- CP-element group 68: 	 branch_block_stmt_1492/if_stmt_1752_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1492/if_stmt_1752_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1492/if_stmt_1752_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1492/if_stmt_1752_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1492/R_cmp_1753_place
      -- CP-element group 68: 	 branch_block_stmt_1492/if_stmt_1752_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1492/if_stmt_1752_else_link/$entry
      -- 
    branch_req_4359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(68), ack => if_stmt_1752_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(52) & convTransposeA_CP_3763_elements(59) & convTransposeA_CP_3763_elements(65) & convTransposeA_CP_3763_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1492/merge_stmt_1758_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/assign_stmt_1764__entry__
      -- CP-element group 69: 	 branch_block_stmt_1492/assign_stmt_1764__exit__
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1492/merge_stmt_1758__exit__
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1492/merge_stmt_1758_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1492/merge_stmt_1758_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1492/merge_stmt_1758_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1492/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/if_stmt_1752_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1492/if_stmt_1752_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1492/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1492/assign_stmt_1764/$entry
      -- CP-element group 69: 	 branch_block_stmt_1492/assign_stmt_1764/$exit
      -- 
    if_choice_transition_4364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1752_branch_ack_1, ack => convTransposeA_CP_3763_elements(69)); -- 
    rr_4704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1822_inst_req_0); -- 
    cr_4709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1822_inst_req_1); -- 
    cr_4732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1816_inst_req_1); -- 
    rr_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1828_inst_req_0); -- 
    cr_4686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1828_inst_req_1); -- 
    rr_4727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1816_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1492/merge_stmt_1766_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1492/merge_stmt_1766__exit__
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802__entry__
      -- CP-element group 70: 	 branch_block_stmt_1492/merge_stmt_1766_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1492/merge_stmt_1766_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1492/merge_stmt_1766_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1492/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1492/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1492/if_stmt_1752_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1492/if_stmt_1752_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1492/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/$entry
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_Update/cr
      -- 
    else_choice_transition_4368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1752_branch_ack_0, ack => convTransposeA_CP_3763_elements(70)); -- 
    rr_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(70), ack => type_cast_1780_inst_req_0); -- 
    cr_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(70), ack => type_cast_1780_inst_req_1); -- 
    cr_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(70), ack => type_cast_1796_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_Sample/ra
      -- 
    ra_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1780_inst_ack_0, ack => convTransposeA_CP_3763_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1780_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_Sample/rr
      -- 
    ca_4390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1780_inst_ack_1, ack => convTransposeA_CP_3763_elements(72)); -- 
    rr_4398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(72), ack => type_cast_1796_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_Sample/ra
      -- 
    ra_4399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1796_inst_ack_0, ack => convTransposeA_CP_3763_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802__exit__
      -- CP-element group 74: 	 branch_block_stmt_1492/if_stmt_1803__entry__
      -- CP-element group 74: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/$exit
      -- CP-element group 74: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1492/assign_stmt_1772_to_assign_stmt_1802/type_cast_1796_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1492/if_stmt_1803_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1492/if_stmt_1803_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1492/if_stmt_1803_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1492/if_stmt_1803_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1492/R_cmp112_1804_place
      -- CP-element group 74: 	 branch_block_stmt_1492/if_stmt_1803_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1492/if_stmt_1803_else_link/$entry
      -- 
    ca_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1796_inst_ack_1, ack => convTransposeA_CP_3763_elements(74)); -- 
    branch_req_4412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(74), ack => if_stmt_1803_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1492/merge_stmt_1837_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1492/merge_stmt_1837_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1492/assign_stmt_1842__entry__
      -- CP-element group 75: 	 branch_block_stmt_1492/merge_stmt_1837__exit__
      -- CP-element group 75: 	 branch_block_stmt_1492/merge_stmt_1837_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1492/merge_stmt_1837_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1492/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1492/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1492/if_stmt_1803_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1492/if_stmt_1803_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1492/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1492/assign_stmt_1842/$entry
      -- CP-element group 75: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_Sample/req
      -- 
    if_choice_transition_4417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1803_branch_ack_1, ack => convTransposeA_CP_3763_elements(75)); -- 
    req_4437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(75), ack => WPIPE_Block0_done_1839_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1810/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1492/if_stmt_1803_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1492/if_stmt_1803_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123
      -- 
    else_choice_transition_4421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1803_branch_ack_0, ack => convTransposeA_CP_3763_elements(76)); -- 
    cr_4629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(76), ack => type_cast_1826_inst_req_1); -- 
    rr_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(76), ack => type_cast_1826_inst_req_0); -- 
    cr_4652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(76), ack => type_cast_1820_inst_req_1); -- 
    rr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(76), ack => type_cast_1820_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_Update/req
      -- 
    ack_4438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1839_inst_ack_0, ack => convTransposeA_CP_3763_elements(77)); -- 
    req_4442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(77), ack => WPIPE_Block0_done_1839_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1492/merge_stmt_1844_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1492/merge_stmt_1844_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1492/merge_stmt_1844_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1492/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1492/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1492/merge_stmt_1844_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1492/assign_stmt_1842__exit__
      -- CP-element group 78: 	 branch_block_stmt_1492/return__
      -- CP-element group 78: 	 branch_block_stmt_1492/branch_block_stmt_1492__exit__
      -- CP-element group 78: 	 branch_block_stmt_1492/merge_stmt_1844__exit__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1492/$exit
      -- CP-element group 78: 	 branch_block_stmt_1492/assign_stmt_1842/$exit
      -- CP-element group 78: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1492/assign_stmt_1842/WPIPE_Block0_done_1839_Update/ack
      -- 
    ack_4443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1839_inst_ack_1, ack => convTransposeA_CP_3763_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1601/$exit
      -- CP-element group 79: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1605_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_req
      -- 
    phi_stmt_1601_req_4454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1601_req_4454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(79), ack => phi_stmt_1601_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(43), ack => convTransposeA_CP_3763_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_req
      -- CP-element group 80: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1612_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1608/$exit
      -- 
    phi_stmt_1608_req_4462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1608_req_4462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(80), ack => phi_stmt_1608_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(43), ack => convTransposeA_CP_3763_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1615/$exit
      -- CP-element group 81: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_req
      -- CP-element group 81: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1619_konst_delay_trans
      -- 
    phi_stmt_1615_req_4470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1615_req_4470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(81), ack => phi_stmt_1615_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(43), ack => convTransposeA_CP_3763_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1622/$exit
      -- CP-element group 82: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1626_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_req
      -- 
    phi_stmt_1622_req_4478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1622_req_4478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(82), ack => phi_stmt_1622_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(43), ack => convTransposeA_CP_3763_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1492/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(79) & convTransposeA_CP_3763_elements(80) & convTransposeA_CP_3763_elements(81) & convTransposeA_CP_3763_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/Sample/ra
      -- 
    ra_4498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_0, ack => convTransposeA_CP_3763_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/Update/ca
      -- 
    ca_4503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_1, ack => convTransposeA_CP_3763_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_req
      -- CP-element group 86: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/type_cast_1607/$exit
      -- CP-element group 86: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/phi_stmt_1601_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1601/$exit
      -- 
    phi_stmt_1601_req_4504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1601_req_4504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(86), ack => phi_stmt_1601_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(84) & convTransposeA_CP_3763_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/Sample/$exit
      -- 
    ra_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1614_inst_ack_0, ack => convTransposeA_CP_3763_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/Update/ca
      -- 
    ca_4526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1614_inst_ack_1, ack => convTransposeA_CP_3763_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_req
      -- CP-element group 89: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/$exit
      -- CP-element group 89: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/type_cast_1614/$exit
      -- CP-element group 89: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1608/phi_stmt_1608_sources/$exit
      -- 
    phi_stmt_1608_req_4527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1608_req_4527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(89), ack => phi_stmt_1608_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(87) & convTransposeA_CP_3763_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/Sample/$exit
      -- 
    ra_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1621_inst_ack_0, ack => convTransposeA_CP_3763_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/Update/$exit
      -- 
    ca_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1621_inst_ack_1, ack => convTransposeA_CP_3763_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_req
      -- CP-element group 92: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/$exit
      -- CP-element group 92: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/$exit
      -- CP-element group 92: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1615/phi_stmt_1615_sources/type_cast_1621/SplitProtocol/$exit
      -- 
    phi_stmt_1615_req_4550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1615_req_4550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(92), ack => phi_stmt_1615_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(90) & convTransposeA_CP_3763_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/Sample/$exit
      -- 
    ra_4567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1628_inst_ack_0, ack => convTransposeA_CP_3763_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/Update/ca
      -- CP-element group 94: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/Update/$exit
      -- 
    ca_4572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1628_inst_ack_1, ack => convTransposeA_CP_3763_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/$exit
      -- CP-element group 95: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_req
      -- CP-element group 95: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1622/phi_stmt_1622_sources/type_cast_1628/$exit
      -- 
    phi_stmt_1622_req_4573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1622_req_4573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(95), ack => phi_stmt_1622_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(93) & convTransposeA_CP_3763_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1492/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(86) & convTransposeA_CP_3763_elements(89) & convTransposeA_CP_3763_elements(92) & convTransposeA_CP_3763_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1492/merge_stmt_1600_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_1492/merge_stmt_1600_PhiAck/$entry
      -- 
    convTransposeA_CP_3763_elements(97) <= OrReduce(convTransposeA_CP_3763_elements(83) & convTransposeA_CP_3763_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1492/merge_stmt_1600_PhiAck/phi_stmt_1601_ack
      -- 
    phi_stmt_1601_ack_4578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1601_ack_0, ack => convTransposeA_CP_3763_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1492/merge_stmt_1600_PhiAck/phi_stmt_1608_ack
      -- 
    phi_stmt_1608_ack_4579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1608_ack_0, ack => convTransposeA_CP_3763_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1492/merge_stmt_1600_PhiAck/phi_stmt_1615_ack
      -- 
    phi_stmt_1615_ack_4580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1615_ack_0, ack => convTransposeA_CP_3763_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1492/merge_stmt_1600_PhiAck/phi_stmt_1622_ack
      -- 
    phi_stmt_1622_ack_4581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1622_ack_0, ack => convTransposeA_CP_3763_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1492/merge_stmt_1600__exit__
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751__entry__
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1663_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1667_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1671_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1701_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1707_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1708_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1712_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/merge_stmt_1600_PhiAck/$exit
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/array_obj_ref_1730_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/addr_of_1731_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/ptr_deref_1734_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1492/assign_stmt_1635_to_assign_stmt_1751/type_cast_1739_Update/cr
      -- 
    rr_4097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1663_inst_req_0); -- 
    cr_4102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1663_inst_req_1); -- 
    rr_4111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1667_inst_req_0); -- 
    cr_4116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1667_inst_req_1); -- 
    rr_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1671_inst_req_0); -- 
    cr_4130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1671_inst_req_1); -- 
    rr_4139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1701_inst_req_0); -- 
    cr_4144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1701_inst_req_1); -- 
    req_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => array_obj_ref_1707_index_offset_req_1); -- 
    req_4190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => addr_of_1708_final_reg_req_1); -- 
    cr_4235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => ptr_deref_1712_load_0_req_1); -- 
    req_4271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => array_obj_ref_1730_index_offset_req_1); -- 
    req_4286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => addr_of_1731_final_reg_req_1); -- 
    cr_4336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => ptr_deref_1734_store_0_req_1); -- 
    rr_4345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1739_inst_req_0); -- 
    cr_4350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(102), ack => type_cast_1739_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(98) & convTransposeA_CP_3763_elements(99) & convTransposeA_CP_3763_elements(100) & convTransposeA_CP_3763_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Sample/$exit
      -- 
    ra_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_0, ack => convTransposeA_CP_3763_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/Update/ca
      -- 
    ca_4630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1826_inst_ack_1, ack => convTransposeA_CP_3763_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	110 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/$exit
      -- CP-element group 105: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/$exit
      -- CP-element group 105: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1826/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_req
      -- 
    phi_stmt_1823_req_4631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1823_req_4631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(105), ack => phi_stmt_1823_req_0); -- 
    convTransposeA_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(103) & convTransposeA_CP_3763_elements(104);
      gj_convTransposeA_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/Sample/ra
      -- 
    ra_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1820_inst_ack_0, ack => convTransposeA_CP_3763_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/Update/ca
      -- CP-element group 107: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/Update/$exit
      -- 
    ca_4653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1820_inst_ack_1, ack => convTransposeA_CP_3763_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/$exit
      -- CP-element group 108: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/$exit
      -- CP-element group 108: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1820/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_req
      -- 
    phi_stmt_1817_req_4654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1817_req_4654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(108), ack => phi_stmt_1817_req_0); -- 
    convTransposeA_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(106) & convTransposeA_CP_3763_elements(107);
      gj_convTransposeA_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  output  delay-element  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_req
      -- CP-element group 109: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1814_konst_delay_trans
      -- CP-element group 109: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1810/$exit
      -- 
    phi_stmt_1810_req_4662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1810_req_4662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(109), ack => phi_stmt_1810_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(76), ack => convTransposeA_CP_3763_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1492/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(105) & convTransposeA_CP_3763_elements(108) & convTransposeA_CP_3763_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Sample/ra
      -- 
    ra_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_0, ack => convTransposeA_CP_3763_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/ca
      -- CP-element group 112: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/Update/$exit
      -- 
    ca_4687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_1, ack => convTransposeA_CP_3763_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/$exit
      -- CP-element group 113: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/$exit
      -- CP-element group 113: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/type_cast_1828/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_sources/$exit
      -- CP-element group 113: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1823/phi_stmt_1823_req
      -- 
    phi_stmt_1823_req_4688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1823_req_4688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(113), ack => phi_stmt_1823_req_1); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(111) & convTransposeA_CP_3763_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/Sample/$exit
      -- 
    ra_4705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1822_inst_ack_0, ack => convTransposeA_CP_3763_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/Update/ca
      -- 
    ca_4710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1822_inst_ack_1, ack => convTransposeA_CP_3763_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_req
      -- CP-element group 116: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/type_cast_1822/$exit
      -- CP-element group 116: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/phi_stmt_1817_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1817/$exit
      -- 
    phi_stmt_1817_req_4711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1817_req_4711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(116), ack => phi_stmt_1817_req_1); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(114) & convTransposeA_CP_3763_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/Sample/ra
      -- 
    ra_4728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1816_inst_ack_0, ack => convTransposeA_CP_3763_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/Update/ca
      -- CP-element group 118: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/Update/$exit
      -- 
    ca_4733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1816_inst_ack_1, ack => convTransposeA_CP_3763_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/$exit
      -- CP-element group 119: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_req
      -- CP-element group 119: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/$exit
      -- CP-element group 119: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1816/SplitProtocol/$exit
      -- 
    phi_stmt_1810_req_4734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1810_req_4734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(119), ack => phi_stmt_1810_req_1); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(117) & convTransposeA_CP_3763_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1492/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(113) & convTransposeA_CP_3763_elements(116) & convTransposeA_CP_3763_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1492/merge_stmt_1809_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_1492/merge_stmt_1809_PhiReqMerge
      -- 
    convTransposeA_CP_3763_elements(121) <= OrReduce(convTransposeA_CP_3763_elements(110) & convTransposeA_CP_3763_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1492/merge_stmt_1809_PhiAck/phi_stmt_1810_ack
      -- 
    phi_stmt_1810_ack_4739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1810_ack_0, ack => convTransposeA_CP_3763_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1492/merge_stmt_1809_PhiAck/phi_stmt_1817_ack
      -- 
    phi_stmt_1817_ack_4740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1817_ack_0, ack => convTransposeA_CP_3763_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1492/merge_stmt_1809_PhiAck/phi_stmt_1823_ack
      -- 
    phi_stmt_1823_ack_4741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1823_ack_0, ack => convTransposeA_CP_3763_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1492/merge_stmt_1809_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(122) & convTransposeA_CP_3763_elements(123) & convTransposeA_CP_3763_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1729_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1729_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1706_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1706_scaled : std_logic_vector(13 downto 0);
    signal add41_1560 : std_logic_vector(15 downto 0);
    signal add54_1571 : std_logic_vector(15 downto 0);
    signal add73_1682 : std_logic_vector(63 downto 0);
    signal add75_1692 : std_logic_vector(63 downto 0);
    signal add86_1746 : std_logic_vector(31 downto 0);
    signal add93_1764 : std_logic_vector(15 downto 0);
    signal add_1544 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1640 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1707_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1707_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1707_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1707_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1707_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1707_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1730_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1730_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1730_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1730_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1730_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1730_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1709 : std_logic_vector(31 downto 0);
    signal arrayidx82_1732 : std_logic_vector(31 downto 0);
    signal call11_1513 : std_logic_vector(15 downto 0);
    signal call13_1516 : std_logic_vector(15 downto 0);
    signal call14_1519 : std_logic_vector(15 downto 0);
    signal call15_1522 : std_logic_vector(15 downto 0);
    signal call16_1535 : std_logic_vector(15 downto 0);
    signal call18_1547 : std_logic_vector(15 downto 0);
    signal call1_1498 : std_logic_vector(15 downto 0);
    signal call20_1550 : std_logic_vector(15 downto 0);
    signal call22_1553 : std_logic_vector(15 downto 0);
    signal call3_1501 : std_logic_vector(15 downto 0);
    signal call5_1504 : std_logic_vector(15 downto 0);
    signal call7_1507 : std_logic_vector(15 downto 0);
    signal call9_1510 : std_logic_vector(15 downto 0);
    signal call_1495 : std_logic_vector(15 downto 0);
    signal cmp101_1777 : std_logic_vector(0 downto 0);
    signal cmp112_1802 : std_logic_vector(0 downto 0);
    signal cmp_1751 : std_logic_vector(0 downto 0);
    signal conv107_1797 : std_logic_vector(31 downto 0);
    signal conv110_1592 : std_logic_vector(31 downto 0);
    signal conv17_1539 : std_logic_vector(31 downto 0);
    signal conv61_1664 : std_logic_vector(63 downto 0);
    signal conv64_1580 : std_logic_vector(63 downto 0);
    signal conv66_1668 : std_logic_vector(63 downto 0);
    signal conv69_1584 : std_logic_vector(63 downto 0);
    signal conv71_1672 : std_logic_vector(63 downto 0);
    signal conv85_1740 : std_logic_vector(31 downto 0);
    signal conv89_1588 : std_logic_vector(31 downto 0);
    signal conv_1526 : std_logic_vector(31 downto 0);
    signal idxprom81_1725 : std_logic_vector(63 downto 0);
    signal idxprom_1702 : std_logic_vector(63 downto 0);
    signal inc105_1781 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1786 : std_logic_vector(15 downto 0);
    signal inc_1772 : std_logic_vector(15 downto 0);
    signal indvar_1601 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1835 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1823 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1622 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1817 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1615 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1793 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1810 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1608 : std_logic_vector(15 downto 0);
    signal mul50_1655 : std_logic_vector(15 downto 0);
    signal mul72_1677 : std_logic_vector(63 downto 0);
    signal mul74_1687 : std_logic_vector(63 downto 0);
    signal mul_1645 : std_logic_vector(15 downto 0);
    signal ptr_deref_1712_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1712_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1712_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1712_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1712_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1734_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1734_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1734_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1734_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1734_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1734_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1532 : std_logic_vector(31 downto 0);
    signal shr111126_1598 : std_logic_vector(31 downto 0);
    signal shr80_1719 : std_logic_vector(63 downto 0);
    signal shr_1698 : std_logic_vector(31 downto 0);
    signal sub44_1650 : std_logic_vector(15 downto 0);
    signal sub57_1576 : std_logic_vector(15 downto 0);
    signal sub58_1660 : std_logic_vector(15 downto 0);
    signal sub_1565 : std_logic_vector(15 downto 0);
    signal tmp1_1635 : std_logic_vector(31 downto 0);
    signal tmp78_1713 : std_logic_vector(63 downto 0);
    signal type_cast_1530_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1558_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1569_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1596_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1605_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1607_wire : std_logic_vector(31 downto 0);
    signal type_cast_1612_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1614_wire : std_logic_vector(15 downto 0);
    signal type_cast_1619_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1621_wire : std_logic_vector(15 downto 0);
    signal type_cast_1626_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1628_wire : std_logic_vector(15 downto 0);
    signal type_cast_1633_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1696_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1717_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1723_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1744_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1762_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1770_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1790_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1814_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1816_wire : std_logic_vector(15 downto 0);
    signal type_cast_1820_wire : std_logic_vector(15 downto 0);
    signal type_cast_1822_wire : std_logic_vector(15 downto 0);
    signal type_cast_1826_wire : std_logic_vector(15 downto 0);
    signal type_cast_1828_wire : std_logic_vector(15 downto 0);
    signal type_cast_1833_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1841_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1707_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1707_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1707_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1707_resized_base_address <= "00000000000000";
    array_obj_ref_1730_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1730_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1730_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1730_resized_base_address <= "00000000000000";
    ptr_deref_1712_word_offset_0 <= "00000000000000";
    ptr_deref_1734_word_offset_0 <= "00000000000000";
    type_cast_1530_wire_constant <= "00000000000000000000000000010000";
    type_cast_1558_wire_constant <= "1111111111111111";
    type_cast_1569_wire_constant <= "1111111111111111";
    type_cast_1596_wire_constant <= "00000000000000000000000000000010";
    type_cast_1605_wire_constant <= "00000000000000000000000000000000";
    type_cast_1612_wire_constant <= "0000000000000000";
    type_cast_1619_wire_constant <= "0000000000000000";
    type_cast_1626_wire_constant <= "0000000000000000";
    type_cast_1633_wire_constant <= "00000000000000000000000000000100";
    type_cast_1696_wire_constant <= "00000000000000000000000000000010";
    type_cast_1717_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1723_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1744_wire_constant <= "00000000000000000000000000000100";
    type_cast_1762_wire_constant <= "0000000000000100";
    type_cast_1770_wire_constant <= "0000000000000001";
    type_cast_1790_wire_constant <= "0000000000000000";
    type_cast_1814_wire_constant <= "0000000000000000";
    type_cast_1833_wire_constant <= "00000000000000000000000000000001";
    type_cast_1841_wire_constant <= "0000000000000001";
    phi_stmt_1601: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1605_wire_constant & type_cast_1607_wire;
      req <= phi_stmt_1601_req_0 & phi_stmt_1601_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1601",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1601_ack_0,
          idata => idata,
          odata => indvar_1601,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1601
    phi_stmt_1608: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1612_wire_constant & type_cast_1614_wire;
      req <= phi_stmt_1608_req_0 & phi_stmt_1608_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1608",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1608_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1608,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1608
    phi_stmt_1615: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1619_wire_constant & type_cast_1621_wire;
      req <= phi_stmt_1615_req_0 & phi_stmt_1615_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1615",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1615_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1615,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1615
    phi_stmt_1622: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1626_wire_constant & type_cast_1628_wire;
      req <= phi_stmt_1622_req_0 & phi_stmt_1622_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1622",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1622_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1622,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1622
    phi_stmt_1810: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1814_wire_constant & type_cast_1816_wire;
      req <= phi_stmt_1810_req_0 & phi_stmt_1810_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1810",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1810_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1810,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1810
    phi_stmt_1817: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1820_wire & type_cast_1822_wire;
      req <= phi_stmt_1817_req_0 & phi_stmt_1817_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1817",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1817_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1817,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1817
    phi_stmt_1823: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1826_wire & type_cast_1828_wire;
      req <= phi_stmt_1823_req_0 & phi_stmt_1823_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1823",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1823_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1823,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1823
    -- flow-through select operator MUX_1792_inst
    input_dim1x_x2_1793 <= type_cast_1790_wire_constant when (cmp101_1777(0) /=  '0') else inc_1772;
    addr_of_1708_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1708_final_reg_req_0;
      addr_of_1708_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1708_final_reg_req_1;
      addr_of_1708_final_reg_ack_1<= rack(0);
      addr_of_1708_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1708_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1707_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1709,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1731_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1731_final_reg_req_0;
      addr_of_1731_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1731_final_reg_req_1;
      addr_of_1731_final_reg_ack_1<= rack(0);
      addr_of_1731_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1731_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1730_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1525_inst_req_0;
      type_cast_1525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1525_inst_req_1;
      type_cast_1525_inst_ack_1<= rack(0);
      type_cast_1525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1522,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1538_inst_req_0;
      type_cast_1538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1538_inst_req_1;
      type_cast_1538_inst_ack_1<= rack(0);
      type_cast_1538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1579_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1579_inst_req_0;
      type_cast_1579_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1579_inst_req_1;
      type_cast_1579_inst_ack_1<= rack(0);
      type_cast_1579_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1579_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1580,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1583_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1583_inst_req_0;
      type_cast_1583_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1583_inst_req_1;
      type_cast_1583_inst_ack_1<= rack(0);
      type_cast_1583_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1583_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1550,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1584,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1587_inst_req_0;
      type_cast_1587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1587_inst_req_1;
      type_cast_1587_inst_ack_1<= rack(0);
      type_cast_1587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1591_inst_req_0;
      type_cast_1591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1591_inst_req_1;
      type_cast_1591_inst_ack_1<= rack(0);
      type_cast_1591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1591_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1592,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1607_inst_req_0;
      type_cast_1607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1607_inst_req_1;
      type_cast_1607_inst_ack_1<= rack(0);
      type_cast_1607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1835,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1607_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1614_inst_req_0;
      type_cast_1614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1614_inst_req_1;
      type_cast_1614_inst_ack_1<= rack(0);
      type_cast_1614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1614_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1621_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1621_inst_req_0;
      type_cast_1621_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1621_inst_req_1;
      type_cast_1621_inst_ack_1<= rack(0);
      type_cast_1621_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1621_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1817,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1621_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1628_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1628_inst_req_0;
      type_cast_1628_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1628_inst_req_1;
      type_cast_1628_inst_ack_1<= rack(0);
      type_cast_1628_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1628_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1823,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1628_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1663_inst_req_0;
      type_cast_1663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1663_inst_req_1;
      type_cast_1663_inst_ack_1<= rack(0);
      type_cast_1663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1663_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1667_inst_req_0;
      type_cast_1667_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1667_inst_req_1;
      type_cast_1667_inst_ack_1<= rack(0);
      type_cast_1667_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1667_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1668,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1671_inst_req_0;
      type_cast_1671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1671_inst_req_1;
      type_cast_1671_inst_ack_1<= rack(0);
      type_cast_1671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1650,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1701_inst_req_0;
      type_cast_1701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1701_inst_req_1;
      type_cast_1701_inst_ack_1<= rack(0);
      type_cast_1701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1739_inst_req_0;
      type_cast_1739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1739_inst_req_1;
      type_cast_1739_inst_ack_1<= rack(0);
      type_cast_1739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1740,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1780_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1780_inst_req_0;
      type_cast_1780_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1780_inst_req_1;
      type_cast_1780_inst_ack_1<= rack(0);
      type_cast_1780_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1780_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1781,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1796_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1796_inst_req_0;
      type_cast_1796_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1796_inst_req_1;
      type_cast_1796_inst_ack_1<= rack(0);
      type_cast_1796_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1796_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1816_inst_req_0;
      type_cast_1816_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1816_inst_req_1;
      type_cast_1816_inst_ack_1<= rack(0);
      type_cast_1816_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1816_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1816_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1820_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1820_inst_req_0;
      type_cast_1820_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1820_inst_req_1;
      type_cast_1820_inst_ack_1<= rack(0);
      type_cast_1820_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1820_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1793,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1820_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1822_inst_req_0;
      type_cast_1822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1822_inst_req_1;
      type_cast_1822_inst_ack_1<= rack(0);
      type_cast_1822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1615,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1822_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1826_inst_req_0;
      type_cast_1826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1826_inst_req_1;
      type_cast_1826_inst_ack_1<= rack(0);
      type_cast_1826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1826_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1828_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1828_inst_req_0;
      type_cast_1828_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1828_inst_req_1;
      type_cast_1828_inst_ack_1<= rack(0);
      type_cast_1828_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1828_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1828_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1707_index_1_rename
    process(R_idxprom_1706_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1706_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1706_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1707_index_1_resize
    process(idxprom_1702) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1702;
      ov := iv(13 downto 0);
      R_idxprom_1706_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1707_root_address_inst
    process(array_obj_ref_1707_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1707_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1707_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1730_index_1_rename
    process(R_idxprom81_1729_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1729_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1729_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1730_index_1_resize
    process(idxprom81_1725) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1725;
      ov := iv(13 downto 0);
      R_idxprom81_1729_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1730_root_address_inst
    process(array_obj_ref_1730_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1730_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1730_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1712_addr_0
    process(ptr_deref_1712_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1712_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1712_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1712_base_resize
    process(arrayidx77_1709) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1709;
      ov := iv(13 downto 0);
      ptr_deref_1712_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1712_gather_scatter
    process(ptr_deref_1712_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1712_data_0;
      ov(63 downto 0) := iv;
      tmp78_1713 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1712_root_address_inst
    process(ptr_deref_1712_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1712_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1712_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1734_addr_0
    process(ptr_deref_1734_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1734_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1734_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1734_base_resize
    process(arrayidx82_1732) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1732;
      ov := iv(13 downto 0);
      ptr_deref_1734_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1734_gather_scatter
    process(tmp78_1713) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1713;
      ov(63 downto 0) := iv;
      ptr_deref_1734_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1734_root_address_inst
    process(ptr_deref_1734_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1734_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1734_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1752_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1751;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1752_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1752_branch_req_0,
          ack0 => if_stmt_1752_branch_ack_0,
          ack1 => if_stmt_1752_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1803_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1802;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1803_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1803_branch_req_0,
          ack0 => if_stmt_1803_branch_ack_0,
          ack1 => if_stmt_1803_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1559_inst
    process(call7_1507) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1507, type_cast_1558_wire_constant, tmp_var);
      add41_1560 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1570_inst
    process(call9_1510) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1510, type_cast_1569_wire_constant, tmp_var);
      add54_1571 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1649_inst
    process(sub_1565, mul_1645) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1565, mul_1645, tmp_var);
      sub44_1650 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1659_inst
    process(sub57_1576, mul50_1655) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1576, mul50_1655, tmp_var);
      sub58_1660 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1763_inst
    process(input_dim2x_x1_1608) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1608, type_cast_1762_wire_constant, tmp_var);
      add93_1764 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1771_inst
    process(input_dim1x_x1_1615) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1615, type_cast_1770_wire_constant, tmp_var);
      inc_1772 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1785_inst
    process(inc105_1781, input_dim0x_x2_1622) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1781, input_dim0x_x2_1622, tmp_var);
      inc105x_xinput_dim0x_x2_1786 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1639_inst
    process(add_1544, tmp1_1635) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1544, tmp1_1635, tmp_var);
      add_src_0x_x0_1640 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1745_inst
    process(conv85_1740) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1740, type_cast_1744_wire_constant, tmp_var);
      add86_1746 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1834_inst
    process(indvar_1601) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1601, type_cast_1833_wire_constant, tmp_var);
      indvarx_xnext_1835 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1681_inst
    process(mul72_1677, conv66_1668) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1677, conv66_1668, tmp_var);
      add73_1682 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1691_inst
    process(mul74_1687, conv61_1664) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1687, conv61_1664, tmp_var);
      add75_1692 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1724_inst
    process(shr80_1719) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1719, type_cast_1723_wire_constant, tmp_var);
      idxprom81_1725 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1776_inst
    process(inc_1772, call1_1498) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1772, call1_1498, tmp_var);
      cmp101_1777 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1801_inst
    process(conv107_1797, shr111126_1598) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1797, shr111126_1598, tmp_var);
      cmp112_1802 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1597_inst
    process(conv110_1592) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1592, type_cast_1596_wire_constant, tmp_var);
      shr111126_1598 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1697_inst
    process(add_src_0x_x0_1640) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1640, type_cast_1696_wire_constant, tmp_var);
      shr_1698 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1718_inst
    process(add75_1692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1692, type_cast_1717_wire_constant, tmp_var);
      shr80_1719 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1644_inst
    process(input_dim0x_x2_1622, call13_1516) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1622, call13_1516, tmp_var);
      mul_1645 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1654_inst
    process(input_dim1x_x1_1615, call13_1516) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1615, call13_1516, tmp_var);
      mul50_1655 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1634_inst
    process(indvar_1601) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1601, type_cast_1633_wire_constant, tmp_var);
      tmp1_1635 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1676_inst
    process(conv71_1672, conv69_1584) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1672, conv69_1584, tmp_var);
      mul72_1677 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1686_inst
    process(add73_1682, conv64_1580) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1682, conv64_1580, tmp_var);
      mul74_1687 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1543_inst
    process(shl_1532, conv17_1539) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1532, conv17_1539, tmp_var);
      add_1544 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1531_inst
    process(conv_1526) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1526, type_cast_1530_wire_constant, tmp_var);
      shl_1532 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1564_inst
    process(add41_1560, call14_1519) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1560, call14_1519, tmp_var);
      sub_1565 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1575_inst
    process(add54_1571, call14_1519) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1571, call14_1519, tmp_var);
      sub57_1576 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1750_inst
    process(add86_1746, conv89_1588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1746, conv89_1588, tmp_var);
      cmp_1751 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1707_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1706_scaled;
      array_obj_ref_1707_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1707_index_offset_req_0;
      array_obj_ref_1707_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1707_index_offset_req_1;
      array_obj_ref_1707_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1730_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1729_scaled;
      array_obj_ref_1730_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1730_index_offset_req_0;
      array_obj_ref_1730_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1730_index_offset_req_1;
      array_obj_ref_1730_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1712_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1712_load_0_req_0;
      ptr_deref_1712_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1712_load_0_req_1;
      ptr_deref_1712_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1712_word_address_0;
      ptr_deref_1712_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1734_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1734_store_0_req_0;
      ptr_deref_1734_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1734_store_0_req_1;
      ptr_deref_1734_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1734_word_address_0;
      data_in <= ptr_deref_1734_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1546_inst RPIPE_Block0_start_1497_inst RPIPE_Block0_start_1500_inst RPIPE_Block0_start_1503_inst RPIPE_Block0_start_1494_inst RPIPE_Block0_start_1549_inst RPIPE_Block0_start_1552_inst RPIPE_Block0_start_1521_inst RPIPE_Block0_start_1518_inst RPIPE_Block0_start_1534_inst RPIPE_Block0_start_1515_inst RPIPE_Block0_start_1512_inst RPIPE_Block0_start_1509_inst RPIPE_Block0_start_1506_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1546_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1497_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1500_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1503_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1494_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1549_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1552_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1521_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1518_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1534_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1515_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1512_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1509_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1506_inst_req_0;
      RPIPE_Block0_start_1546_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1497_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1500_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1503_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1494_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1549_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1552_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1521_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1518_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1534_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1515_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1512_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1509_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1506_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1546_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1497_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1500_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1503_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1494_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1549_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1552_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1521_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1518_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1534_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1515_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1512_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1509_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1506_inst_req_1;
      RPIPE_Block0_start_1546_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1497_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1500_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1503_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1494_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1549_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1552_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1521_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1518_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1534_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1515_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1512_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1509_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1506_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call18_1547 <= data_out(223 downto 208);
      call1_1498 <= data_out(207 downto 192);
      call3_1501 <= data_out(191 downto 176);
      call5_1504 <= data_out(175 downto 160);
      call_1495 <= data_out(159 downto 144);
      call20_1550 <= data_out(143 downto 128);
      call22_1553 <= data_out(127 downto 112);
      call15_1522 <= data_out(111 downto 96);
      call14_1519 <= data_out(95 downto 80);
      call16_1535 <= data_out(79 downto 64);
      call13_1516 <= data_out(63 downto 48);
      call11_1513 <= data_out(47 downto 32);
      call9_1510 <= data_out(31 downto 16);
      call7_1507 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1839_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1839_inst_req_0;
      WPIPE_Block0_done_1839_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1839_inst_req_1;
      WPIPE_Block0_done_1839_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1841_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4758_start: Boolean;
  signal convTransposeB_CP_4758_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1868_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1874_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1859_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1865_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1877_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1868_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1868_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1877_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1865_inst_ack_1 : boolean;
  signal type_cast_1894_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1877_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1902_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1859_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1859_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1874_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1850_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1865_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1865_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1862_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1850_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1853_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1853_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1850_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1859_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1905_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1902_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1902_inst_req_1 : boolean;
  signal type_cast_1945_inst_req_0 : boolean;
  signal type_cast_1945_inst_ack_0 : boolean;
  signal type_cast_1894_inst_ack_1 : boolean;
  signal type_cast_1894_inst_req_1 : boolean;
  signal type_cast_1941_inst_req_1 : boolean;
  signal type_cast_1941_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1908_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1908_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1902_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1877_inst_req_1 : boolean;
  signal type_cast_1881_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1874_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1874_inst_req_1 : boolean;
  signal type_cast_1881_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1850_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1868_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1905_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1856_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1905_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1856_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1905_inst_req_1 : boolean;
  signal type_cast_1894_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1890_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1890_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1871_inst_ack_1 : boolean;
  signal type_cast_1953_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1871_inst_req_1 : boolean;
  signal type_cast_1953_inst_req_0 : boolean;
  signal type_cast_1953_inst_ack_0 : boolean;
  signal type_cast_1953_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1890_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1890_inst_req_0 : boolean;
  signal type_cast_2024_inst_req_1 : boolean;
  signal type_cast_2024_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1871_inst_ack_0 : boolean;
  signal type_cast_1945_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1871_inst_req_0 : boolean;
  signal type_cast_1949_inst_req_0 : boolean;
  signal type_cast_1949_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1853_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1862_inst_ack_1 : boolean;
  signal type_cast_1949_inst_req_1 : boolean;
  signal type_cast_1949_inst_ack_1 : boolean;
  signal type_cast_2181_inst_req_0 : boolean;
  signal type_cast_2024_inst_req_0 : boolean;
  signal type_cast_2024_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1853_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1862_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1856_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1856_inst_req_0 : boolean;
  signal type_cast_1945_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1862_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1908_inst_req_1 : boolean;
  signal type_cast_1881_inst_ack_0 : boolean;
  signal type_cast_1941_inst_req_0 : boolean;
  signal type_cast_1941_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1908_inst_ack_1 : boolean;
  signal type_cast_1881_inst_req_0 : boolean;
  signal phi_stmt_2171_req_1 : boolean;
  signal type_cast_2028_inst_req_0 : boolean;
  signal type_cast_2028_inst_ack_0 : boolean;
  signal type_cast_2028_inst_req_1 : boolean;
  signal type_cast_2028_inst_ack_1 : boolean;
  signal phi_stmt_2171_req_0 : boolean;
  signal type_cast_2032_inst_req_0 : boolean;
  signal type_cast_2032_inst_ack_0 : boolean;
  signal type_cast_2183_inst_req_1 : boolean;
  signal type_cast_2032_inst_req_1 : boolean;
  signal type_cast_2032_inst_ack_1 : boolean;
  signal type_cast_2174_inst_ack_1 : boolean;
  signal type_cast_2062_inst_req_0 : boolean;
  signal type_cast_2062_inst_ack_0 : boolean;
  signal type_cast_2062_inst_req_1 : boolean;
  signal type_cast_2062_inst_ack_1 : boolean;
  signal type_cast_2174_inst_req_1 : boolean;
  signal type_cast_2174_inst_ack_0 : boolean;
  signal type_cast_2174_inst_req_0 : boolean;
  signal array_obj_ref_2068_index_offset_req_0 : boolean;
  signal array_obj_ref_2068_index_offset_ack_0 : boolean;
  signal array_obj_ref_2068_index_offset_req_1 : boolean;
  signal array_obj_ref_2068_index_offset_ack_1 : boolean;
  signal addr_of_2069_final_reg_req_0 : boolean;
  signal addr_of_2069_final_reg_ack_0 : boolean;
  signal addr_of_2069_final_reg_req_1 : boolean;
  signal addr_of_2069_final_reg_ack_1 : boolean;
  signal type_cast_2187_inst_ack_0 : boolean;
  signal type_cast_2187_inst_req_0 : boolean;
  signal ptr_deref_2073_load_0_req_0 : boolean;
  signal ptr_deref_2073_load_0_ack_0 : boolean;
  signal ptr_deref_2073_load_0_req_1 : boolean;
  signal ptr_deref_2073_load_0_ack_1 : boolean;
  signal type_cast_2183_inst_ack_0 : boolean;
  signal phi_stmt_2184_req_1 : boolean;
  signal array_obj_ref_2091_index_offset_req_0 : boolean;
  signal array_obj_ref_2091_index_offset_ack_0 : boolean;
  signal array_obj_ref_2091_index_offset_req_1 : boolean;
  signal array_obj_ref_2091_index_offset_ack_1 : boolean;
  signal type_cast_2189_inst_ack_1 : boolean;
  signal addr_of_2092_final_reg_req_0 : boolean;
  signal addr_of_2092_final_reg_ack_0 : boolean;
  signal addr_of_2092_final_reg_req_1 : boolean;
  signal addr_of_2092_final_reg_ack_1 : boolean;
  signal type_cast_2189_inst_req_1 : boolean;
  signal type_cast_2183_inst_req_0 : boolean;
  signal ptr_deref_2095_store_0_req_0 : boolean;
  signal type_cast_2189_inst_ack_0 : boolean;
  signal ptr_deref_2095_store_0_ack_0 : boolean;
  signal ptr_deref_2095_store_0_req_1 : boolean;
  signal ptr_deref_2095_store_0_ack_1 : boolean;
  signal type_cast_2189_inst_req_0 : boolean;
  signal type_cast_2100_inst_req_0 : boolean;
  signal type_cast_2100_inst_ack_0 : boolean;
  signal type_cast_2100_inst_req_1 : boolean;
  signal type_cast_2100_inst_ack_1 : boolean;
  signal if_stmt_2113_branch_req_0 : boolean;
  signal if_stmt_2113_branch_ack_1 : boolean;
  signal phi_stmt_2184_ack_0 : boolean;
  signal if_stmt_2113_branch_ack_0 : boolean;
  signal phi_stmt_2178_ack_0 : boolean;
  signal phi_stmt_2171_ack_0 : boolean;
  signal type_cast_2141_inst_req_0 : boolean;
  signal type_cast_2141_inst_ack_0 : boolean;
  signal type_cast_2141_inst_req_1 : boolean;
  signal type_cast_2141_inst_ack_1 : boolean;
  signal type_cast_2157_inst_req_0 : boolean;
  signal type_cast_2157_inst_ack_0 : boolean;
  signal type_cast_2157_inst_req_1 : boolean;
  signal type_cast_2157_inst_ack_1 : boolean;
  signal phi_stmt_2178_req_0 : boolean;
  signal if_stmt_2164_branch_req_0 : boolean;
  signal type_cast_2181_inst_ack_1 : boolean;
  signal if_stmt_2164_branch_ack_1 : boolean;
  signal type_cast_2181_inst_req_1 : boolean;
  signal if_stmt_2164_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2200_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2200_inst_ack_0 : boolean;
  signal phi_stmt_2184_req_0 : boolean;
  signal WPIPE_Block1_done_2200_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2200_inst_ack_1 : boolean;
  signal type_cast_1987_inst_req_0 : boolean;
  signal type_cast_1987_inst_ack_0 : boolean;
  signal type_cast_1987_inst_req_1 : boolean;
  signal type_cast_1987_inst_ack_1 : boolean;
  signal phi_stmt_1984_req_0 : boolean;
  signal type_cast_2187_inst_ack_1 : boolean;
  signal phi_stmt_1977_req_0 : boolean;
  signal phi_stmt_1970_req_0 : boolean;
  signal phi_stmt_1963_req_1 : boolean;
  signal type_cast_1989_inst_req_0 : boolean;
  signal type_cast_1989_inst_ack_0 : boolean;
  signal type_cast_1989_inst_req_1 : boolean;
  signal type_cast_1989_inst_ack_1 : boolean;
  signal phi_stmt_1984_req_1 : boolean;
  signal type_cast_2187_inst_req_1 : boolean;
  signal type_cast_1983_inst_req_0 : boolean;
  signal type_cast_1983_inst_ack_0 : boolean;
  signal type_cast_1983_inst_req_1 : boolean;
  signal type_cast_1983_inst_ack_1 : boolean;
  signal phi_stmt_1977_req_1 : boolean;
  signal type_cast_1976_inst_req_0 : boolean;
  signal type_cast_1976_inst_ack_0 : boolean;
  signal type_cast_1976_inst_req_1 : boolean;
  signal type_cast_1976_inst_ack_1 : boolean;
  signal phi_stmt_1970_req_1 : boolean;
  signal type_cast_1966_inst_req_0 : boolean;
  signal type_cast_1966_inst_ack_0 : boolean;
  signal type_cast_1966_inst_req_1 : boolean;
  signal phi_stmt_2178_req_1 : boolean;
  signal type_cast_1966_inst_ack_1 : boolean;
  signal phi_stmt_1963_req_0 : boolean;
  signal type_cast_2181_inst_ack_0 : boolean;
  signal type_cast_2183_inst_ack_1 : boolean;
  signal phi_stmt_1963_ack_0 : boolean;
  signal phi_stmt_1970_ack_0 : boolean;
  signal phi_stmt_1977_ack_0 : boolean;
  signal phi_stmt_1984_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4758_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4758_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4758_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4758_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4758: Block -- control-path 
    signal convTransposeB_CP_4758_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4758_elements(0) <= convTransposeB_CP_4758_start;
    convTransposeB_CP_4758_symbol <= convTransposeB_CP_4758_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909__entry__
      -- CP-element group 0: 	 branch_block_stmt_1848/branch_block_stmt_1848__entry__
      -- CP-element group 0: 	 branch_block_stmt_1848/$entry
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/$entry
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_update_start_
      -- 
    rr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(0), ack => RPIPE_Block1_start_1850_inst_req_0); -- 
    cr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(0), ack => type_cast_1894_inst_req_1); -- 
    cr_4951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(0), ack => type_cast_1881_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1848/assign_stmt_2196__entry__
      -- CP-element group 1: 	 branch_block_stmt_1848/assign_stmt_2196__exit__
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1848/merge_stmt_2170__exit__
      -- CP-element group 1: 	 branch_block_stmt_1848/assign_stmt_2196/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/assign_stmt_2196/$exit
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/Update/cr
      -- 
    rr_5507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1989_inst_req_0); -- 
    cr_5512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1989_inst_req_1); -- 
    rr_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1983_inst_req_0); -- 
    cr_5535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1983_inst_req_1); -- 
    rr_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1976_inst_req_0); -- 
    cr_5558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1976_inst_req_1); -- 
    rr_5576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1966_inst_req_0); -- 
    cr_5581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(1), ack => type_cast_1966_inst_req_1); -- 
    convTransposeB_CP_4758_elements(1) <= convTransposeB_CP_4758_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_Update/cr
      -- 
    ra_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1850_inst_ack_0, ack => convTransposeB_CP_4758_elements(2)); -- 
    cr_4811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(2), ack => RPIPE_Block1_start_1850_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1850_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_Sample/$entry
      -- 
    ca_4812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1850_inst_ack_1, ack => convTransposeB_CP_4758_elements(3)); -- 
    rr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(3), ack => RPIPE_Block1_start_1853_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_update_start_
      -- 
    ra_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1853_inst_ack_0, ack => convTransposeB_CP_4758_elements(4)); -- 
    cr_4825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(4), ack => RPIPE_Block1_start_1853_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1853_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_sample_start_
      -- 
    ca_4826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1853_inst_ack_1, ack => convTransposeB_CP_4758_elements(5)); -- 
    rr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(5), ack => RPIPE_Block1_start_1856_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_Sample/$exit
      -- 
    ra_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1856_inst_ack_0, ack => convTransposeB_CP_4758_elements(6)); -- 
    cr_4839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(6), ack => RPIPE_Block1_start_1856_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1856_Update/$exit
      -- 
    ca_4840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1856_inst_ack_1, ack => convTransposeB_CP_4758_elements(7)); -- 
    rr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(7), ack => RPIPE_Block1_start_1859_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_sample_completed_
      -- 
    ra_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1859_inst_ack_0, ack => convTransposeB_CP_4758_elements(8)); -- 
    cr_4853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(8), ack => RPIPE_Block1_start_1859_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1859_Update/$exit
      -- 
    ca_4854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1859_inst_ack_1, ack => convTransposeB_CP_4758_elements(9)); -- 
    rr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(9), ack => RPIPE_Block1_start_1862_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_Sample/ra
      -- 
    ra_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1862_inst_ack_0, ack => convTransposeB_CP_4758_elements(10)); -- 
    cr_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(10), ack => RPIPE_Block1_start_1862_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1862_Update/$exit
      -- 
    ca_4868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1862_inst_ack_1, ack => convTransposeB_CP_4758_elements(11)); -- 
    rr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(11), ack => RPIPE_Block1_start_1865_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_sample_completed_
      -- 
    ra_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1865_inst_ack_0, ack => convTransposeB_CP_4758_elements(12)); -- 
    cr_4881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(12), ack => RPIPE_Block1_start_1865_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1865_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_Sample/$entry
      -- 
    ca_4882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1865_inst_ack_1, ack => convTransposeB_CP_4758_elements(13)); -- 
    rr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(13), ack => RPIPE_Block1_start_1868_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_Sample/$exit
      -- 
    ra_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1868_inst_ack_0, ack => convTransposeB_CP_4758_elements(14)); -- 
    cr_4895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(14), ack => RPIPE_Block1_start_1868_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1868_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_Sample/$entry
      -- 
    ca_4896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1868_inst_ack_1, ack => convTransposeB_CP_4758_elements(15)); -- 
    rr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(15), ack => RPIPE_Block1_start_1871_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_update_start_
      -- 
    ra_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1871_inst_ack_0, ack => convTransposeB_CP_4758_elements(16)); -- 
    cr_4909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(16), ack => RPIPE_Block1_start_1871_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1871_Update/$exit
      -- 
    ca_4910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1871_inst_ack_1, ack => convTransposeB_CP_4758_elements(17)); -- 
    rr_4918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(17), ack => RPIPE_Block1_start_1874_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_sample_completed_
      -- 
    ra_4919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1874_inst_ack_0, ack => convTransposeB_CP_4758_elements(18)); -- 
    cr_4923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(18), ack => RPIPE_Block1_start_1874_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1874_update_completed_
      -- 
    ca_4924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1874_inst_ack_1, ack => convTransposeB_CP_4758_elements(19)); -- 
    rr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(19), ack => RPIPE_Block1_start_1877_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_Update/$entry
      -- 
    ra_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1877_inst_ack_0, ack => convTransposeB_CP_4758_elements(20)); -- 
    cr_4937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(20), ack => RPIPE_Block1_start_1877_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1877_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_Sample/$entry
      -- 
    ca_4938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1877_inst_ack_1, ack => convTransposeB_CP_4758_elements(21)); -- 
    rr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(21), ack => type_cast_1881_inst_req_0); -- 
    rr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(21), ack => RPIPE_Block1_start_1890_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_Sample/$exit
      -- 
    ra_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_0, ack => convTransposeB_CP_4758_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1881_Update/$exit
      -- 
    ca_4952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_1, ack => convTransposeB_CP_4758_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_sample_completed_
      -- 
    ra_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1890_inst_ack_0, ack => convTransposeB_CP_4758_elements(24)); -- 
    cr_4965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(24), ack => RPIPE_Block1_start_1890_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1890_update_completed_
      -- 
    ca_4966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1890_inst_ack_1, ack => convTransposeB_CP_4758_elements(25)); -- 
    rr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(25), ack => type_cast_1894_inst_req_0); -- 
    rr_4988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(25), ack => RPIPE_Block1_start_1902_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_sample_completed_
      -- 
    ra_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1894_inst_ack_0, ack => convTransposeB_CP_4758_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/type_cast_1894_update_completed_
      -- 
    ca_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1894_inst_ack_1, ack => convTransposeB_CP_4758_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_update_start_
      -- 
    ra_4989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1902_inst_ack_0, ack => convTransposeB_CP_4758_elements(28)); -- 
    cr_4993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(28), ack => RPIPE_Block1_start_1902_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1902_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_Sample/rr
      -- 
    ca_4994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1902_inst_ack_1, ack => convTransposeB_CP_4758_elements(29)); -- 
    rr_5002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(29), ack => RPIPE_Block1_start_1905_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_Update/cr
      -- 
    ra_5003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1905_inst_ack_0, ack => convTransposeB_CP_4758_elements(30)); -- 
    cr_5007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(30), ack => RPIPE_Block1_start_1905_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1905_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_Sample/$entry
      -- 
    ca_5008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1905_inst_ack_1, ack => convTransposeB_CP_4758_elements(31)); -- 
    rr_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(31), ack => RPIPE_Block1_start_1908_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_Update/cr
      -- 
    ra_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1908_inst_ack_0, ack => convTransposeB_CP_4758_elements(32)); -- 
    cr_5021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(32), ack => RPIPE_Block1_start_1908_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/RPIPE_Block1_start_1908_Update/ca
      -- 
    ca_5022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1908_inst_ack_1, ack => convTransposeB_CP_4758_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909__exit__
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960__entry__
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1851_to_assign_stmt_1909/$exit
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_update_start_
      -- 
    rr_5047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1945_inst_req_0); -- 
    cr_5038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1941_inst_req_1); -- 
    cr_5080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1953_inst_req_1); -- 
    rr_5075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1953_inst_req_0); -- 
    cr_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1945_inst_req_1); -- 
    rr_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1949_inst_req_0); -- 
    cr_5066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1949_inst_req_1); -- 
    rr_5033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(34), ack => type_cast_1941_inst_req_0); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(23) & convTransposeB_CP_4758_elements(27) & convTransposeB_CP_4758_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_Sample/ra
      -- 
    ra_5034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_0, ack => convTransposeB_CP_4758_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1941_update_completed_
      -- 
    ca_5039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_1, ack => convTransposeB_CP_4758_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_Sample/$exit
      -- 
    ra_5048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_0, ack => convTransposeB_CP_4758_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1945_Update/ca
      -- 
    ca_5053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_1, ack => convTransposeB_CP_4758_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_sample_completed_
      -- 
    ra_5062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1949_inst_ack_0, ack => convTransposeB_CP_4758_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1949_update_completed_
      -- 
    ca_5067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1949_inst_ack_1, ack => convTransposeB_CP_4758_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_sample_completed_
      -- 
    ra_5076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_0, ack => convTransposeB_CP_4758_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/type_cast_1953_update_completed_
      -- 
    ca_5081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_1, ack => convTransposeB_CP_4758_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960__exit__
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1848/assign_stmt_1916_to_assign_stmt_1960/$exit
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1977/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1970/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1963/$entry
      -- CP-element group 43: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/$entry
      -- 
    rr_5457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(43), ack => type_cast_1987_inst_req_0); -- 
    cr_5462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(43), ack => type_cast_1987_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(36) & convTransposeB_CP_4758_elements(38) & convTransposeB_CP_4758_elements(40) & convTransposeB_CP_4758_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_Sample/ra
      -- 
    ra_5093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2024_inst_ack_0, ack => convTransposeB_CP_4758_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_Update/$exit
      -- 
    ca_5098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2024_inst_ack_1, ack => convTransposeB_CP_4758_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_Sample/ra
      -- 
    ra_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2028_inst_ack_0, ack => convTransposeB_CP_4758_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_Update/ca
      -- 
    ca_5112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2028_inst_ack_1, ack => convTransposeB_CP_4758_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_Sample/ra
      -- 
    ra_5121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2032_inst_ack_0, ack => convTransposeB_CP_4758_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_Update/ca
      -- 
    ca_5126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2032_inst_ack_1, ack => convTransposeB_CP_4758_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_Sample/ra
      -- 
    ra_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2062_inst_ack_0, ack => convTransposeB_CP_4758_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_Sample/req
      -- 
    ca_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2062_inst_ack_1, ack => convTransposeB_CP_4758_elements(51)); -- 
    req_5165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(51), ack => array_obj_ref_2068_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_Sample/ack
      -- 
    ack_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2068_index_offset_ack_0, ack => convTransposeB_CP_4758_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_request/req
      -- 
    ack_5171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2068_index_offset_ack_1, ack => convTransposeB_CP_4758_elements(53)); -- 
    req_5180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(53), ack => addr_of_2069_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_request/ack
      -- 
    ack_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2069_final_reg_ack_0, ack => convTransposeB_CP_4758_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Sample/word_access_start/word_0/rr
      -- 
    ack_5186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2069_final_reg_ack_1, ack => convTransposeB_CP_4758_elements(55)); -- 
    rr_5219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(55), ack => ptr_deref_2073_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Sample/word_access_start/word_0/ra
      -- 
    ra_5220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2073_load_0_ack_0, ack => convTransposeB_CP_4758_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/ptr_deref_2073_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/ptr_deref_2073_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/ptr_deref_2073_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/ptr_deref_2073_Merge/merge_ack
      -- 
    ca_5231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2073_load_0_ack_1, ack => convTransposeB_CP_4758_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_Sample/req
      -- 
    req_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(58), ack => array_obj_ref_2091_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(45) & convTransposeB_CP_4758_elements(47) & convTransposeB_CP_4758_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_Sample/ack
      -- 
    ack_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2091_index_offset_ack_0, ack => convTransposeB_CP_4758_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_request/req
      -- 
    ack_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2091_index_offset_ack_1, ack => convTransposeB_CP_4758_elements(60)); -- 
    req_5276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(60), ack => addr_of_2092_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_request/ack
      -- 
    ack_5277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2092_final_reg_ack_0, ack => convTransposeB_CP_4758_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_word_addrgen/root_register_ack
      -- 
    ack_5282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2092_final_reg_ack_1, ack => convTransposeB_CP_4758_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/ptr_deref_2095_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/ptr_deref_2095_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/ptr_deref_2095_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/ptr_deref_2095_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/word_access_start/word_0/rr
      -- 
    rr_5320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(63), ack => ptr_deref_2095_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(57) & convTransposeB_CP_4758_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Sample/word_access_start/word_0/ra
      -- 
    ra_5321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2095_store_0_ack_0, ack => convTransposeB_CP_4758_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Update/word_access_complete/word_0/ca
      -- 
    ca_5332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2095_store_0_ack_1, ack => convTransposeB_CP_4758_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_Sample/ra
      -- 
    ra_5341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2100_inst_ack_0, ack => convTransposeB_CP_4758_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_Update/ca
      -- 
    ca_5346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2100_inst_ack_1, ack => convTransposeB_CP_4758_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112__exit__
      -- CP-element group 68: 	 branch_block_stmt_1848/if_stmt_2113__entry__
      -- CP-element group 68: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/$exit
      -- CP-element group 68: 	 branch_block_stmt_1848/if_stmt_2113_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1848/if_stmt_2113_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1848/if_stmt_2113_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1848/if_stmt_2113_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1848/R_cmp_2114_place
      -- CP-element group 68: 	 branch_block_stmt_1848/if_stmt_2113_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1848/if_stmt_2113_else_link/$entry
      -- 
    branch_req_5354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(68), ack => if_stmt_2113_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(52) & convTransposeB_CP_4758_elements(59) & convTransposeB_CP_4758_elements(65) & convTransposeB_CP_4758_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1848/merge_stmt_2119__exit__
      -- CP-element group 69: 	 branch_block_stmt_1848/assign_stmt_2125__entry__
      -- CP-element group 69: 	 branch_block_stmt_1848/assign_stmt_2125__exit__
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1848/if_stmt_2113_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1848/if_stmt_2113_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1848/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1848/assign_stmt_2125/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/assign_stmt_2125/$exit
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/merge_stmt_2119_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/merge_stmt_2119_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/merge_stmt_2119_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1848/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1848/merge_stmt_2119_PhiReqMerge
      -- 
    if_choice_transition_5359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2113_branch_ack_1, ack => convTransposeB_CP_4758_elements(69)); -- 
    rr_5737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2181_inst_req_0); -- 
    cr_5719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2174_inst_req_1); -- 
    rr_5714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2174_inst_req_0); -- 
    cr_5696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2189_inst_req_1); -- 
    rr_5691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2189_inst_req_0); -- 
    cr_5742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(69), ack => type_cast_2181_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1848/merge_stmt_2127__exit__
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163__entry__
      -- CP-element group 70: 	 branch_block_stmt_1848/merge_stmt_2127_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1848/merge_stmt_2127_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1848/merge_stmt_2127_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1848/if_stmt_2113_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1848/if_stmt_2113_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1848/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/$entry
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1848/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1848/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1848/merge_stmt_2127_PhiReqMerge
      -- 
    else_choice_transition_5363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2113_branch_ack_0, ack => convTransposeB_CP_4758_elements(70)); -- 
    rr_5379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(70), ack => type_cast_2141_inst_req_0); -- 
    cr_5384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(70), ack => type_cast_2141_inst_req_1); -- 
    cr_5398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(70), ack => type_cast_2157_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_Sample/ra
      -- 
    ra_5380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2141_inst_ack_0, ack => convTransposeB_CP_4758_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2141_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_Sample/rr
      -- 
    ca_5385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2141_inst_ack_1, ack => convTransposeB_CP_4758_elements(72)); -- 
    rr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(72), ack => type_cast_2157_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_Sample/ra
      -- 
    ra_5394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2157_inst_ack_0, ack => convTransposeB_CP_4758_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163__exit__
      -- CP-element group 74: 	 branch_block_stmt_1848/if_stmt_2164__entry__
      -- CP-element group 74: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/$exit
      -- CP-element group 74: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1848/assign_stmt_2133_to_assign_stmt_2163/type_cast_2157_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1848/if_stmt_2164_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1848/if_stmt_2164_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1848/if_stmt_2164_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1848/if_stmt_2164_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1848/R_cmp117_2165_place
      -- CP-element group 74: 	 branch_block_stmt_1848/if_stmt_2164_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1848/if_stmt_2164_else_link/$entry
      -- 
    ca_5399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2157_inst_ack_1, ack => convTransposeB_CP_4758_elements(74)); -- 
    branch_req_5407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(74), ack => if_stmt_2164_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1848/assign_stmt_2203__entry__
      -- CP-element group 75: 	 branch_block_stmt_1848/merge_stmt_2198__exit__
      -- CP-element group 75: 	 branch_block_stmt_1848/merge_stmt_2198_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1848/merge_stmt_2198_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1848/merge_stmt_2198_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1848/merge_stmt_2198_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1848/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1848/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1848/if_stmt_2164_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1848/if_stmt_2164_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1848/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1848/assign_stmt_2203/$entry
      -- CP-element group 75: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_Sample/req
      -- 
    if_choice_transition_5412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2164_branch_ack_1, ack => convTransposeB_CP_4758_elements(75)); -- 
    req_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(75), ack => WPIPE_Block1_done_2200_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	108 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2171/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/if_stmt_2164_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1848/if_stmt_2164_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/$entry
      -- 
    else_choice_transition_5416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2164_branch_ack_0, ack => convTransposeB_CP_4758_elements(76)); -- 
    cr_5670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(76), ack => type_cast_2183_inst_req_1); -- 
    rr_5634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(76), ack => type_cast_2187_inst_req_0); -- 
    rr_5665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(76), ack => type_cast_2183_inst_req_0); -- 
    cr_5639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(76), ack => type_cast_2187_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_Update/req
      -- 
    ack_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2200_inst_ack_0, ack => convTransposeB_CP_4758_elements(77)); -- 
    req_5437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(77), ack => WPIPE_Block1_done_2200_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1848/branch_block_stmt_1848__exit__
      -- CP-element group 78: 	 branch_block_stmt_1848/$exit
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1848/merge_stmt_2205__exit__
      -- CP-element group 78: 	 branch_block_stmt_1848/return__
      -- CP-element group 78: 	 branch_block_stmt_1848/assign_stmt_2203__exit__
      -- CP-element group 78: 	 branch_block_stmt_1848/merge_stmt_2205_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1848/merge_stmt_2205_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1848/merge_stmt_2205_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1848/merge_stmt_2205_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1848/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1848/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1848/assign_stmt_2203/$exit
      -- CP-element group 78: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1848/assign_stmt_2203/WPIPE_Block1_done_2200_Update/ack
      -- 
    ack_5438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2200_inst_ack_1, ack => convTransposeB_CP_4758_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Sample/ra
      -- 
    ra_5458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1987_inst_ack_0, ack => convTransposeB_CP_4758_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/Update/ca
      -- 
    ca_5463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1987_inst_ack_1, ack => convTransposeB_CP_4758_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/$exit
      -- CP-element group 81: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/$exit
      -- CP-element group 81: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1987/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_req
      -- 
    phi_stmt_1984_req_5464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1984_req_5464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(81), ack => phi_stmt_1984_req_0); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(79) & convTransposeB_CP_4758_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1977/$exit
      -- CP-element group 82: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1981_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_req
      -- 
    phi_stmt_1977_req_5472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1977_req_5472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(82), ack => phi_stmt_1977_req_0); -- 
    -- Element group convTransposeB_CP_4758_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4758_elements(43), ack => convTransposeB_CP_4758_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1970/$exit
      -- CP-element group 83: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1974_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_req
      -- 
    phi_stmt_1970_req_5480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1970_req_5480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(83), ack => phi_stmt_1970_req_0); -- 
    -- Element group convTransposeB_CP_4758_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4758_elements(43), ack => convTransposeB_CP_4758_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1963/$exit
      -- CP-element group 84: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1969_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_req
      -- 
    phi_stmt_1963_req_5488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1963_req_5488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(84), ack => phi_stmt_1963_req_1); -- 
    -- Element group convTransposeB_CP_4758_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4758_elements(43), ack => convTransposeB_CP_4758_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1848/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(81) & convTransposeB_CP_4758_elements(82) & convTransposeB_CP_4758_elements(83) & convTransposeB_CP_4758_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Sample/ra
      -- 
    ra_5508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1989_inst_ack_0, ack => convTransposeB_CP_4758_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/Update/ca
      -- 
    ca_5513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1989_inst_ack_1, ack => convTransposeB_CP_4758_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/$exit
      -- CP-element group 88: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/$exit
      -- CP-element group 88: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_sources/type_cast_1989/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1984/phi_stmt_1984_req
      -- 
    phi_stmt_1984_req_5514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1984_req_5514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(88), ack => phi_stmt_1984_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(86) & convTransposeB_CP_4758_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/Sample/ra
      -- 
    ra_5531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1983_inst_ack_0, ack => convTransposeB_CP_4758_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/Update/ca
      -- 
    ca_5536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1983_inst_ack_1, ack => convTransposeB_CP_4758_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/$exit
      -- CP-element group 91: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/$exit
      -- CP-element group 91: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_sources/type_cast_1983/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1977/phi_stmt_1977_req
      -- 
    phi_stmt_1977_req_5537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1977_req_5537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(91), ack => phi_stmt_1977_req_1); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(89) & convTransposeB_CP_4758_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/Sample/ra
      -- 
    ra_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_0, ack => convTransposeB_CP_4758_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/Update/ca
      -- 
    ca_5559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_1, ack => convTransposeB_CP_4758_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/$exit
      -- CP-element group 94: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/$exit
      -- CP-element group 94: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_sources/type_cast_1976/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1970/phi_stmt_1970_req
      -- 
    phi_stmt_1970_req_5560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1970_req_5560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(94), ack => phi_stmt_1970_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(92) & convTransposeB_CP_4758_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/Sample/ra
      -- 
    ra_5577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1966_inst_ack_0, ack => convTransposeB_CP_4758_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/Update/ca
      -- 
    ca_5582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1966_inst_ack_1, ack => convTransposeB_CP_4758_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/$exit
      -- CP-element group 97: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/$exit
      -- CP-element group 97: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_sources/type_cast_1966/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1963/phi_stmt_1963_req
      -- 
    phi_stmt_1963_req_5583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1963_req_5583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(97), ack => phi_stmt_1963_req_0); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(95) & convTransposeB_CP_4758_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1848/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(88) & convTransposeB_CP_4758_elements(91) & convTransposeB_CP_4758_elements(94) & convTransposeB_CP_4758_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1848/merge_stmt_1962_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_1848/merge_stmt_1962_PhiAck/$entry
      -- 
    convTransposeB_CP_4758_elements(99) <= OrReduce(convTransposeB_CP_4758_elements(85) & convTransposeB_CP_4758_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1848/merge_stmt_1962_PhiAck/phi_stmt_1963_ack
      -- 
    phi_stmt_1963_ack_5588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1963_ack_0, ack => convTransposeB_CP_4758_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1848/merge_stmt_1962_PhiAck/phi_stmt_1970_ack
      -- 
    phi_stmt_1970_ack_5589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1970_ack_0, ack => convTransposeB_CP_4758_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1848/merge_stmt_1962_PhiAck/phi_stmt_1977_ack
      -- 
    phi_stmt_1977_ack_5590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1977_ack_0, ack => convTransposeB_CP_4758_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1848/merge_stmt_1962_PhiAck/phi_stmt_1984_ack
      -- 
    phi_stmt_1984_ack_5591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1984_ack_0, ack => convTransposeB_CP_4758_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112__entry__
      -- CP-element group 104: 	 branch_block_stmt_1848/merge_stmt_1962__exit__
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2024_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2028_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2032_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2062_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2068_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2069_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2073_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/array_obj_ref_2091_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/addr_of_2092_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/ptr_deref_2095_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1848/assign_stmt_1996_to_assign_stmt_2112/type_cast_2100_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1848/merge_stmt_1962_PhiAck/$exit
      -- 
    cr_5097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2024_inst_req_1); -- 
    rr_5092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2024_inst_req_0); -- 
    rr_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2028_inst_req_0); -- 
    cr_5111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2028_inst_req_1); -- 
    rr_5120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2032_inst_req_0); -- 
    cr_5125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2032_inst_req_1); -- 
    rr_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2062_inst_req_0); -- 
    cr_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2062_inst_req_1); -- 
    req_5170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => array_obj_ref_2068_index_offset_req_1); -- 
    req_5185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => addr_of_2069_final_reg_req_1); -- 
    cr_5230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => ptr_deref_2073_load_0_req_1); -- 
    req_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => array_obj_ref_2091_index_offset_req_1); -- 
    req_5281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => addr_of_2092_final_reg_req_1); -- 
    cr_5331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => ptr_deref_2095_store_0_req_1); -- 
    rr_5340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2100_inst_req_0); -- 
    cr_5345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(104), ack => type_cast_2100_inst_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(100) & convTransposeB_CP_4758_elements(101) & convTransposeB_CP_4758_elements(102) & convTransposeB_CP_4758_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Sample/$exit
      -- 
    ra_5635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_0, ack => convTransposeB_CP_4758_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/Update/ca
      -- 
    ca_5640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2187_inst_ack_1, ack => convTransposeB_CP_4758_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2187/$exit
      -- CP-element group 107: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/$exit
      -- CP-element group 107: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_req
      -- 
    phi_stmt_2184_req_5641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2184_req_5641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(107), ack => phi_stmt_2184_req_0); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(105) & convTransposeB_CP_4758_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  output  delay-element  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2177_konst_delay_trans
      -- CP-element group 108: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_req
      -- CP-element group 108: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2171/$exit
      -- 
    phi_stmt_2171_req_5649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2171_req_5649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(108), ack => phi_stmt_2171_req_1); -- 
    -- Element group convTransposeB_CP_4758_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => convTransposeB_CP_4758_elements(76), ack => convTransposeB_CP_4758_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/Sample/$exit
      -- 
    ra_5666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2183_inst_ack_0, ack => convTransposeB_CP_4758_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/Update/ca
      -- 
    ca_5671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2183_inst_ack_1, ack => convTransposeB_CP_4758_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2183/$exit
      -- CP-element group 111: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/$exit
      -- CP-element group 111: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_req
      -- 
    phi_stmt_2178_req_5672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2178_req_5672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(111), ack => phi_stmt_2178_req_1); -- 
    convTransposeB_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(109) & convTransposeB_CP_4758_elements(110);
      gj_convTransposeB_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1848/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(107) & convTransposeB_CP_4758_elements(108) & convTransposeB_CP_4758_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Sample/$exit
      -- 
    ra_5692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_0, ack => convTransposeB_CP_4758_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Update/ca
      -- CP-element group 114: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/Update/$exit
      -- 
    ca_5697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_1, ack => convTransposeB_CP_4758_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_req
      -- CP-element group 115: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/type_cast_2189/$exit
      -- CP-element group 115: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/phi_stmt_2184_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2184/$exit
      -- 
    phi_stmt_2184_req_5698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2184_req_5698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(115), ack => phi_stmt_2184_req_1); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(113) & convTransposeB_CP_4758_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Sample/$exit
      -- 
    ra_5715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2174_inst_ack_0, ack => convTransposeB_CP_4758_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/Update/$exit
      -- 
    ca_5720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2174_inst_ack_1, ack => convTransposeB_CP_4758_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_req
      -- CP-element group 118: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/type_cast_2174/$exit
      -- CP-element group 118: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/phi_stmt_2171_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2171/$exit
      -- 
    phi_stmt_2171_req_5721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2171_req_5721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(118), ack => phi_stmt_2171_req_0); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(116) & convTransposeB_CP_4758_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/Sample/ra
      -- 
    ra_5738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2181_inst_ack_0, ack => convTransposeB_CP_4758_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/Update/$exit
      -- 
    ca_5743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2181_inst_ack_1, ack => convTransposeB_CP_4758_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/$exit
      -- CP-element group 121: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_sources/type_cast_2181/$exit
      -- CP-element group 121: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2178/phi_stmt_2178_req
      -- 
    phi_stmt_2178_req_5744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2178_req_5744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4758_elements(121), ack => phi_stmt_2178_req_0); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(119) & convTransposeB_CP_4758_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1848/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(115) & convTransposeB_CP_4758_elements(118) & convTransposeB_CP_4758_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1848/merge_stmt_2170_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_1848/merge_stmt_2170_PhiAck/$entry
      -- 
    convTransposeB_CP_4758_elements(123) <= OrReduce(convTransposeB_CP_4758_elements(112) & convTransposeB_CP_4758_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1848/merge_stmt_2170_PhiAck/phi_stmt_2171_ack
      -- 
    phi_stmt_2171_ack_5749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2171_ack_0, ack => convTransposeB_CP_4758_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1848/merge_stmt_2170_PhiAck/phi_stmt_2178_ack
      -- 
    phi_stmt_2178_ack_5750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2178_ack_0, ack => convTransposeB_CP_4758_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1848/merge_stmt_2170_PhiAck/phi_stmt_2184_ack
      -- 
    phi_stmt_2184_ack_5751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2184_ack_0, ack => convTransposeB_CP_4758_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1848/merge_stmt_2170_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4758_elements(124) & convTransposeB_CP_4758_elements(125) & convTransposeB_CP_4758_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4758_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2090_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2090_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2067_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2067_scaled : std_logic_vector(13 downto 0);
    signal add45_1922 : std_logic_vector(15 downto 0);
    signal add58_1933 : std_logic_vector(15 downto 0);
    signal add77_2043 : std_logic_vector(63 downto 0);
    signal add79_2053 : std_logic_vector(63 downto 0);
    signal add91_2107 : std_logic_vector(31 downto 0);
    signal add98_2125 : std_logic_vector(15 downto 0);
    signal add_1900 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2001 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2068_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2068_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2068_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2068_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2068_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2068_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2091_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2091_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2091_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2091_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2091_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2091_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2070 : std_logic_vector(31 downto 0);
    signal arrayidx87_2093 : std_logic_vector(31 downto 0);
    signal call11_1869 : std_logic_vector(15 downto 0);
    signal call13_1872 : std_logic_vector(15 downto 0);
    signal call14_1875 : std_logic_vector(15 downto 0);
    signal call15_1878 : std_logic_vector(15 downto 0);
    signal call16_1891 : std_logic_vector(15 downto 0);
    signal call18_1903 : std_logic_vector(15 downto 0);
    signal call1_1854 : std_logic_vector(15 downto 0);
    signal call20_1906 : std_logic_vector(15 downto 0);
    signal call22_1909 : std_logic_vector(15 downto 0);
    signal call3_1857 : std_logic_vector(15 downto 0);
    signal call5_1860 : std_logic_vector(15 downto 0);
    signal call7_1863 : std_logic_vector(15 downto 0);
    signal call9_1866 : std_logic_vector(15 downto 0);
    signal call_1851 : std_logic_vector(15 downto 0);
    signal cmp106_2138 : std_logic_vector(0 downto 0);
    signal cmp117_2163 : std_logic_vector(0 downto 0);
    signal cmp_2112 : std_logic_vector(0 downto 0);
    signal conv112_2158 : std_logic_vector(31 downto 0);
    signal conv115_1954 : std_logic_vector(31 downto 0);
    signal conv17_1895 : std_logic_vector(31 downto 0);
    signal conv65_2025 : std_logic_vector(63 downto 0);
    signal conv68_1942 : std_logic_vector(63 downto 0);
    signal conv70_2029 : std_logic_vector(63 downto 0);
    signal conv73_1946 : std_logic_vector(63 downto 0);
    signal conv75_2033 : std_logic_vector(63 downto 0);
    signal conv90_2101 : std_logic_vector(31 downto 0);
    signal conv94_1950 : std_logic_vector(31 downto 0);
    signal conv_1882 : std_logic_vector(31 downto 0);
    signal idxprom86_2086 : std_logic_vector(63 downto 0);
    signal idxprom_2063 : std_logic_vector(63 downto 0);
    signal inc110_2142 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2147 : std_logic_vector(15 downto 0);
    signal inc_2133 : std_logic_vector(15 downto 0);
    signal indvar_1963 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2196 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2184 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1984 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2178 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1977 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2154 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2171 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1970 : std_logic_vector(15 downto 0);
    signal mul54_2016 : std_logic_vector(15 downto 0);
    signal mul76_2038 : std_logic_vector(63 downto 0);
    signal mul78_2048 : std_logic_vector(63 downto 0);
    signal mul_2006 : std_logic_vector(15 downto 0);
    signal ptr_deref_2073_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2073_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2073_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2073_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2073_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2095_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2095_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2095_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2095_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2095_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2095_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1888 : std_logic_vector(31 downto 0);
    signal shr116132_1960 : std_logic_vector(31 downto 0);
    signal shr131_1916 : std_logic_vector(15 downto 0);
    signal shr81_2059 : std_logic_vector(31 downto 0);
    signal shr85_2080 : std_logic_vector(63 downto 0);
    signal sub48_2011 : std_logic_vector(15 downto 0);
    signal sub61_1938 : std_logic_vector(15 downto 0);
    signal sub62_2021 : std_logic_vector(15 downto 0);
    signal sub_1927 : std_logic_vector(15 downto 0);
    signal tmp1_1996 : std_logic_vector(31 downto 0);
    signal tmp83_2074 : std_logic_vector(63 downto 0);
    signal type_cast_1886_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1914_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1920_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1931_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1958_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1966_wire : std_logic_vector(31 downto 0);
    signal type_cast_1969_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1974_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1976_wire : std_logic_vector(15 downto 0);
    signal type_cast_1981_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1983_wire : std_logic_vector(15 downto 0);
    signal type_cast_1987_wire : std_logic_vector(15 downto 0);
    signal type_cast_1989_wire : std_logic_vector(15 downto 0);
    signal type_cast_1994_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2057_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2078_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2084_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2105_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2123_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2131_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2151_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2174_wire : std_logic_vector(15 downto 0);
    signal type_cast_2177_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2181_wire : std_logic_vector(15 downto 0);
    signal type_cast_2183_wire : std_logic_vector(15 downto 0);
    signal type_cast_2187_wire : std_logic_vector(15 downto 0);
    signal type_cast_2189_wire : std_logic_vector(15 downto 0);
    signal type_cast_2194_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2202_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2068_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2068_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2068_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2068_resized_base_address <= "00000000000000";
    array_obj_ref_2091_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2091_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2091_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2091_resized_base_address <= "00000000000000";
    ptr_deref_2073_word_offset_0 <= "00000000000000";
    ptr_deref_2095_word_offset_0 <= "00000000000000";
    type_cast_1886_wire_constant <= "00000000000000000000000000010000";
    type_cast_1914_wire_constant <= "0000000000000010";
    type_cast_1920_wire_constant <= "1111111111111111";
    type_cast_1931_wire_constant <= "1111111111111111";
    type_cast_1958_wire_constant <= "00000000000000000000000000000001";
    type_cast_1969_wire_constant <= "00000000000000000000000000000000";
    type_cast_1974_wire_constant <= "0000000000000000";
    type_cast_1981_wire_constant <= "0000000000000000";
    type_cast_1994_wire_constant <= "00000000000000000000000000000100";
    type_cast_2057_wire_constant <= "00000000000000000000000000000010";
    type_cast_2078_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2084_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2105_wire_constant <= "00000000000000000000000000000100";
    type_cast_2123_wire_constant <= "0000000000000100";
    type_cast_2131_wire_constant <= "0000000000000001";
    type_cast_2151_wire_constant <= "0000000000000000";
    type_cast_2177_wire_constant <= "0000000000000000";
    type_cast_2194_wire_constant <= "00000000000000000000000000000001";
    type_cast_2202_wire_constant <= "0000000000000001";
    phi_stmt_1963: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1966_wire & type_cast_1969_wire_constant;
      req <= phi_stmt_1963_req_0 & phi_stmt_1963_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1963",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1963_ack_0,
          idata => idata,
          odata => indvar_1963,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1963
    phi_stmt_1970: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1974_wire_constant & type_cast_1976_wire;
      req <= phi_stmt_1970_req_0 & phi_stmt_1970_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1970",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1970_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1970,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1970
    phi_stmt_1977: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1981_wire_constant & type_cast_1983_wire;
      req <= phi_stmt_1977_req_0 & phi_stmt_1977_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1977",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1977_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1977,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1977
    phi_stmt_1984: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1987_wire & type_cast_1989_wire;
      req <= phi_stmt_1984_req_0 & phi_stmt_1984_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1984",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1984_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1984,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1984
    phi_stmt_2171: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2174_wire & type_cast_2177_wire_constant;
      req <= phi_stmt_2171_req_0 & phi_stmt_2171_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2171",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2171_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2171,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2171
    phi_stmt_2178: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2181_wire & type_cast_2183_wire;
      req <= phi_stmt_2178_req_0 & phi_stmt_2178_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2178",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2178_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2178,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2178
    phi_stmt_2184: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2187_wire & type_cast_2189_wire;
      req <= phi_stmt_2184_req_0 & phi_stmt_2184_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2184",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2184_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2184,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2184
    -- flow-through select operator MUX_2153_inst
    input_dim1x_x2_2154 <= type_cast_2151_wire_constant when (cmp106_2138(0) /=  '0') else inc_2133;
    addr_of_2069_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2069_final_reg_req_0;
      addr_of_2069_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2069_final_reg_req_1;
      addr_of_2069_final_reg_ack_1<= rack(0);
      addr_of_2069_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2069_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2068_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2070,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2092_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2092_final_reg_req_0;
      addr_of_2092_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2092_final_reg_req_1;
      addr_of_2092_final_reg_ack_1<= rack(0);
      addr_of_2092_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2092_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2091_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2093,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1881_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1881_inst_req_0;
      type_cast_1881_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1881_inst_req_1;
      type_cast_1881_inst_ack_1<= rack(0);
      type_cast_1881_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1881_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1878,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1882,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1894_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1894_inst_req_0;
      type_cast_1894_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1894_inst_req_1;
      type_cast_1894_inst_ack_1<= rack(0);
      type_cast_1894_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1894_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1891,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1895,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1941_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1941_inst_req_0;
      type_cast_1941_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1941_inst_req_1;
      type_cast_1941_inst_ack_1<= rack(0);
      type_cast_1941_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1941_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1909,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1942,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1945_inst_req_0;
      type_cast_1945_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1945_inst_req_1;
      type_cast_1945_inst_ack_1<= rack(0);
      type_cast_1945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1906,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1946,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1949_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1949_inst_req_0;
      type_cast_1949_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1949_inst_req_1;
      type_cast_1949_inst_ack_1<= rack(0);
      type_cast_1949_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1949_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1857,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1950,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1953_inst_req_0;
      type_cast_1953_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1953_inst_req_1;
      type_cast_1953_inst_ack_1<= rack(0);
      type_cast_1953_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1953_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1851,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1954,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1966_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1966_inst_req_0;
      type_cast_1966_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1966_inst_req_1;
      type_cast_1966_inst_ack_1<= rack(0);
      type_cast_1966_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1966_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1966_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1976_inst_req_0;
      type_cast_1976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1976_inst_req_1;
      type_cast_1976_inst_ack_1<= rack(0);
      type_cast_1976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1976_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1983_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1983_inst_req_0;
      type_cast_1983_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1983_inst_req_1;
      type_cast_1983_inst_ack_1<= rack(0);
      type_cast_1983_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1983_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2178,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1983_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1987_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1987_inst_req_0;
      type_cast_1987_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1987_inst_req_1;
      type_cast_1987_inst_ack_1<= rack(0);
      type_cast_1987_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1987_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1916,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1987_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1989_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1989_inst_req_0;
      type_cast_1989_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1989_inst_req_1;
      type_cast_1989_inst_ack_1<= rack(0);
      type_cast_1989_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1989_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1989_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2024_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2024_inst_req_0;
      type_cast_2024_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2024_inst_req_1;
      type_cast_2024_inst_ack_1<= rack(0);
      type_cast_2024_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2024_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1970,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2025,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2028_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2028_inst_req_0;
      type_cast_2028_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2028_inst_req_1;
      type_cast_2028_inst_ack_1<= rack(0);
      type_cast_2028_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2028_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2021,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2029,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2032_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2032_inst_req_0;
      type_cast_2032_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2032_inst_req_1;
      type_cast_2032_inst_ack_1<= rack(0);
      type_cast_2032_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2032_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2011,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2033,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2062_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2062_inst_req_0;
      type_cast_2062_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2062_inst_req_1;
      type_cast_2062_inst_ack_1<= rack(0);
      type_cast_2062_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2062_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2059,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2063,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2100_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2100_inst_req_0;
      type_cast_2100_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2100_inst_req_1;
      type_cast_2100_inst_ack_1<= rack(0);
      type_cast_2100_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2100_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1970,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2101,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2141_inst_req_0;
      type_cast_2141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2141_inst_req_1;
      type_cast_2141_inst_ack_1<= rack(0);
      type_cast_2141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2157_inst_req_0;
      type_cast_2157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2157_inst_req_1;
      type_cast_2157_inst_ack_1<= rack(0);
      type_cast_2157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2147,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2174_inst_req_0;
      type_cast_2174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2174_inst_req_1;
      type_cast_2174_inst_ack_1<= rack(0);
      type_cast_2174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2174_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2181_inst_req_0;
      type_cast_2181_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2181_inst_req_1;
      type_cast_2181_inst_ack_1<= rack(0);
      type_cast_2181_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2181_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1977,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2181_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2183_inst_req_0;
      type_cast_2183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2183_inst_req_1;
      type_cast_2183_inst_ack_1<= rack(0);
      type_cast_2183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2183_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2183_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2187_inst_req_0;
      type_cast_2187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2187_inst_req_1;
      type_cast_2187_inst_ack_1<= rack(0);
      type_cast_2187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2147,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2187_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2189_inst_req_0;
      type_cast_2189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2189_inst_req_1;
      type_cast_2189_inst_ack_1<= rack(0);
      type_cast_2189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2189_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2068_index_1_rename
    process(R_idxprom_2067_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2067_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2067_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2068_index_1_resize
    process(idxprom_2063) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2063;
      ov := iv(13 downto 0);
      R_idxprom_2067_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2068_root_address_inst
    process(array_obj_ref_2068_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2068_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2068_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2091_index_1_rename
    process(R_idxprom86_2090_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2090_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2090_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2091_index_1_resize
    process(idxprom86_2086) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2086;
      ov := iv(13 downto 0);
      R_idxprom86_2090_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2091_root_address_inst
    process(array_obj_ref_2091_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2091_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2091_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_addr_0
    process(ptr_deref_2073_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2073_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2073_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_base_resize
    process(arrayidx82_2070) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2070;
      ov := iv(13 downto 0);
      ptr_deref_2073_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_gather_scatter
    process(ptr_deref_2073_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2073_data_0;
      ov(63 downto 0) := iv;
      tmp83_2074 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_root_address_inst
    process(ptr_deref_2073_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2073_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2073_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2095_addr_0
    process(ptr_deref_2095_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2095_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2095_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2095_base_resize
    process(arrayidx87_2093) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2093;
      ov := iv(13 downto 0);
      ptr_deref_2095_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2095_gather_scatter
    process(tmp83_2074) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2074;
      ov(63 downto 0) := iv;
      ptr_deref_2095_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2095_root_address_inst
    process(ptr_deref_2095_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2095_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2095_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2113_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2112;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2113_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2113_branch_req_0,
          ack0 => if_stmt_2113_branch_ack_0,
          ack1 => if_stmt_2113_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2164_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2163;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2164_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2164_branch_req_0,
          ack0 => if_stmt_2164_branch_ack_0,
          ack1 => if_stmt_2164_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1921_inst
    process(call7_1863) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1863, type_cast_1920_wire_constant, tmp_var);
      add45_1922 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1932_inst
    process(call9_1866) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1866, type_cast_1931_wire_constant, tmp_var);
      add58_1933 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2010_inst
    process(sub_1927, mul_2006) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1927, mul_2006, tmp_var);
      sub48_2011 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2020_inst
    process(sub61_1938, mul54_2016) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1938, mul54_2016, tmp_var);
      sub62_2021 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2124_inst
    process(input_dim2x_x1_1970) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1970, type_cast_2123_wire_constant, tmp_var);
      add98_2125 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2132_inst
    process(input_dim1x_x1_1977) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1977, type_cast_2131_wire_constant, tmp_var);
      inc_2133 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2146_inst
    process(inc110_2142, input_dim0x_x2_1984) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2142, input_dim0x_x2_1984, tmp_var);
      inc110x_xinput_dim0x_x2_2147 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2000_inst
    process(add_1900, tmp1_1996) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1900, tmp1_1996, tmp_var);
      add_src_0x_x0_2001 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2106_inst
    process(conv90_2101) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2101, type_cast_2105_wire_constant, tmp_var);
      add91_2107 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2195_inst
    process(indvar_1963) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1963, type_cast_2194_wire_constant, tmp_var);
      indvarx_xnext_2196 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2042_inst
    process(mul76_2038, conv70_2029) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2038, conv70_2029, tmp_var);
      add77_2043 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2052_inst
    process(mul78_2048, conv65_2025) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2048, conv65_2025, tmp_var);
      add79_2053 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2085_inst
    process(shr85_2080) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2080, type_cast_2084_wire_constant, tmp_var);
      idxprom86_2086 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2137_inst
    process(inc_2133, call1_1854) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2133, call1_1854, tmp_var);
      cmp106_2138 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2162_inst
    process(conv112_2158, shr116132_1960) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2158, shr116132_1960, tmp_var);
      cmp117_2163 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1915_inst
    process(call_1851) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1851, type_cast_1914_wire_constant, tmp_var);
      shr131_1916 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1959_inst
    process(conv115_1954) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1954, type_cast_1958_wire_constant, tmp_var);
      shr116132_1960 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2058_inst
    process(add_src_0x_x0_2001) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2001, type_cast_2057_wire_constant, tmp_var);
      shr81_2059 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2079_inst
    process(add79_2053) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2053, type_cast_2078_wire_constant, tmp_var);
      shr85_2080 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2005_inst
    process(input_dim0x_x2_1984, call13_1872) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1984, call13_1872, tmp_var);
      mul_2006 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2015_inst
    process(input_dim1x_x1_1977, call13_1872) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1977, call13_1872, tmp_var);
      mul54_2016 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1995_inst
    process(indvar_1963) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1963, type_cast_1994_wire_constant, tmp_var);
      tmp1_1996 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2037_inst
    process(conv75_2033, conv73_1946) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2033, conv73_1946, tmp_var);
      mul76_2038 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2047_inst
    process(add77_2043, conv68_1942) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2043, conv68_1942, tmp_var);
      mul78_2048 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1899_inst
    process(shl_1888, conv17_1895) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1888, conv17_1895, tmp_var);
      add_1900 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1887_inst
    process(conv_1882) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1882, type_cast_1886_wire_constant, tmp_var);
      shl_1888 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1926_inst
    process(add45_1922, call14_1875) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1922, call14_1875, tmp_var);
      sub_1927 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1937_inst
    process(add58_1933, call14_1875) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1933, call14_1875, tmp_var);
      sub61_1938 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2111_inst
    process(add91_2107, conv94_1950) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2107, conv94_1950, tmp_var);
      cmp_2112 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2068_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2067_scaled;
      array_obj_ref_2068_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2068_index_offset_req_0;
      array_obj_ref_2068_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2068_index_offset_req_1;
      array_obj_ref_2068_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2091_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2090_scaled;
      array_obj_ref_2091_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2091_index_offset_req_0;
      array_obj_ref_2091_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2091_index_offset_req_1;
      array_obj_ref_2091_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_2073_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2073_load_0_req_0;
      ptr_deref_2073_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2073_load_0_req_1;
      ptr_deref_2073_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2073_word_address_0;
      ptr_deref_2073_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2095_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2095_store_0_req_0;
      ptr_deref_2095_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2095_store_0_req_1;
      ptr_deref_2095_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2095_word_address_0;
      data_in <= ptr_deref_2095_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1856_inst RPIPE_Block1_start_1859_inst RPIPE_Block1_start_1865_inst RPIPE_Block1_start_1862_inst RPIPE_Block1_start_1853_inst RPIPE_Block1_start_1850_inst RPIPE_Block1_start_1908_inst RPIPE_Block1_start_1905_inst RPIPE_Block1_start_1902_inst RPIPE_Block1_start_1890_inst RPIPE_Block1_start_1877_inst RPIPE_Block1_start_1874_inst RPIPE_Block1_start_1871_inst RPIPE_Block1_start_1868_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1856_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1859_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1865_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1862_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1853_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1850_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1908_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1905_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1902_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1890_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1877_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1874_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1871_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1868_inst_req_0;
      RPIPE_Block1_start_1856_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1859_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1865_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1862_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1853_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1850_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1908_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1905_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1902_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1890_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1877_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1874_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1871_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1868_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1856_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1859_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1865_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1862_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1853_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1850_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1908_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1905_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1902_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1890_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1877_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1874_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1871_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1868_inst_req_1;
      RPIPE_Block1_start_1856_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1859_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1865_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1862_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1853_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1850_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1908_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1905_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1902_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1890_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1877_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1874_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1871_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1868_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call3_1857 <= data_out(223 downto 208);
      call5_1860 <= data_out(207 downto 192);
      call9_1866 <= data_out(191 downto 176);
      call7_1863 <= data_out(175 downto 160);
      call1_1854 <= data_out(159 downto 144);
      call_1851 <= data_out(143 downto 128);
      call22_1909 <= data_out(127 downto 112);
      call20_1906 <= data_out(111 downto 96);
      call18_1903 <= data_out(95 downto 80);
      call16_1891 <= data_out(79 downto 64);
      call15_1878 <= data_out(63 downto 48);
      call14_1875 <= data_out(47 downto 32);
      call13_1872 <= data_out(31 downto 16);
      call11_1869 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2200_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2200_inst_req_0;
      WPIPE_Block1_done_2200_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2200_inst_req_1;
      WPIPE_Block1_done_2200_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2202_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5768_start: Boolean;
  signal convTransposeC_CP_5768_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block2_start_2232_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2238_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2229_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2266_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2226_inst_ack_0 : boolean;
  signal type_cast_2255_inst_ack_1 : boolean;
  signal type_cast_2242_inst_req_1 : boolean;
  signal type_cast_2242_inst_ack_0 : boolean;
  signal type_cast_2242_inst_ack_1 : boolean;
  signal type_cast_2242_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2263_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2235_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2269_inst_ack_0 : boolean;
  signal type_cast_2255_inst_req_1 : boolean;
  signal type_cast_2306_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2223_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2238_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2263_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2223_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2266_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2251_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2226_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2251_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2251_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2226_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2226_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2238_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2269_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2251_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2238_inst_ack_1 : boolean;
  signal type_cast_2255_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2263_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2269_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2266_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2269_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2263_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2235_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2235_inst_req_1 : boolean;
  signal type_cast_2310_inst_ack_0 : boolean;
  signal type_cast_2310_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2232_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2229_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2229_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2235_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2266_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2229_inst_ack_0 : boolean;
  signal type_cast_2255_inst_req_0 : boolean;
  signal type_cast_2396_inst_ack_0 : boolean;
  signal type_cast_2310_inst_req_0 : boolean;
  signal type_cast_2396_inst_req_0 : boolean;
  signal type_cast_2302_inst_ack_1 : boolean;
  signal type_cast_2302_inst_req_1 : boolean;
  signal type_cast_2314_inst_req_1 : boolean;
  signal type_cast_2314_inst_ack_1 : boolean;
  signal type_cast_2314_inst_req_0 : boolean;
  signal type_cast_2314_inst_ack_0 : boolean;
  signal type_cast_2396_inst_req_1 : boolean;
  signal type_cast_2396_inst_ack_1 : boolean;
  signal type_cast_2306_inst_ack_1 : boolean;
  signal type_cast_2302_inst_ack_0 : boolean;
  signal type_cast_2306_inst_req_1 : boolean;
  signal type_cast_2302_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2232_inst_ack_1 : boolean;
  signal type_cast_2310_inst_req_1 : boolean;
  signal type_cast_2306_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2232_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2223_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2220_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2223_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2220_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2211_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2211_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2211_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2211_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2214_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2214_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2214_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2214_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2217_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2217_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2217_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2217_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2220_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2220_inst_ack_0 : boolean;
  signal type_cast_2400_inst_req_0 : boolean;
  signal type_cast_2400_inst_ack_0 : boolean;
  signal type_cast_2400_inst_req_1 : boolean;
  signal type_cast_2400_inst_ack_1 : boolean;
  signal type_cast_2404_inst_req_0 : boolean;
  signal type_cast_2404_inst_ack_0 : boolean;
  signal type_cast_2404_inst_req_1 : boolean;
  signal type_cast_2404_inst_ack_1 : boolean;
  signal type_cast_2434_inst_req_0 : boolean;
  signal type_cast_2434_inst_ack_0 : boolean;
  signal type_cast_2434_inst_req_1 : boolean;
  signal type_cast_2434_inst_ack_1 : boolean;
  signal array_obj_ref_2440_index_offset_req_0 : boolean;
  signal array_obj_ref_2440_index_offset_ack_0 : boolean;
  signal array_obj_ref_2440_index_offset_req_1 : boolean;
  signal array_obj_ref_2440_index_offset_ack_1 : boolean;
  signal addr_of_2441_final_reg_req_0 : boolean;
  signal addr_of_2441_final_reg_ack_0 : boolean;
  signal addr_of_2441_final_reg_req_1 : boolean;
  signal addr_of_2441_final_reg_ack_1 : boolean;
  signal ptr_deref_2445_load_0_req_0 : boolean;
  signal ptr_deref_2445_load_0_ack_0 : boolean;
  signal ptr_deref_2445_load_0_req_1 : boolean;
  signal ptr_deref_2445_load_0_ack_1 : boolean;
  signal array_obj_ref_2463_index_offset_req_0 : boolean;
  signal array_obj_ref_2463_index_offset_ack_0 : boolean;
  signal array_obj_ref_2463_index_offset_req_1 : boolean;
  signal array_obj_ref_2463_index_offset_ack_1 : boolean;
  signal addr_of_2464_final_reg_req_0 : boolean;
  signal addr_of_2464_final_reg_ack_0 : boolean;
  signal addr_of_2464_final_reg_req_1 : boolean;
  signal addr_of_2464_final_reg_ack_1 : boolean;
  signal ptr_deref_2467_store_0_req_0 : boolean;
  signal ptr_deref_2467_store_0_ack_0 : boolean;
  signal ptr_deref_2467_store_0_req_1 : boolean;
  signal ptr_deref_2467_store_0_ack_1 : boolean;
  signal type_cast_2472_inst_req_0 : boolean;
  signal type_cast_2472_inst_ack_0 : boolean;
  signal type_cast_2472_inst_req_1 : boolean;
  signal type_cast_2472_inst_ack_1 : boolean;
  signal if_stmt_2485_branch_req_0 : boolean;
  signal if_stmt_2485_branch_ack_1 : boolean;
  signal if_stmt_2485_branch_ack_0 : boolean;
  signal type_cast_2513_inst_req_0 : boolean;
  signal type_cast_2513_inst_ack_0 : boolean;
  signal type_cast_2513_inst_req_1 : boolean;
  signal type_cast_2513_inst_ack_1 : boolean;
  signal type_cast_2529_inst_req_0 : boolean;
  signal type_cast_2529_inst_ack_0 : boolean;
  signal type_cast_2529_inst_req_1 : boolean;
  signal type_cast_2529_inst_ack_1 : boolean;
  signal if_stmt_2536_branch_req_0 : boolean;
  signal if_stmt_2536_branch_ack_1 : boolean;
  signal if_stmt_2536_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2572_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2572_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2572_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2572_inst_ack_1 : boolean;
  signal phi_stmt_2335_req_0 : boolean;
  signal phi_stmt_2342_req_0 : boolean;
  signal phi_stmt_2349_req_1 : boolean;
  signal type_cast_2361_inst_req_0 : boolean;
  signal type_cast_2361_inst_ack_0 : boolean;
  signal type_cast_2361_inst_req_1 : boolean;
  signal type_cast_2361_inst_ack_1 : boolean;
  signal phi_stmt_2356_req_1 : boolean;
  signal type_cast_2341_inst_req_0 : boolean;
  signal type_cast_2341_inst_ack_0 : boolean;
  signal type_cast_2341_inst_req_1 : boolean;
  signal type_cast_2341_inst_ack_1 : boolean;
  signal phi_stmt_2335_req_1 : boolean;
  signal type_cast_2348_inst_req_0 : boolean;
  signal type_cast_2348_inst_ack_0 : boolean;
  signal type_cast_2348_inst_req_1 : boolean;
  signal type_cast_2348_inst_ack_1 : boolean;
  signal phi_stmt_2342_req_1 : boolean;
  signal type_cast_2352_inst_req_0 : boolean;
  signal type_cast_2352_inst_ack_0 : boolean;
  signal type_cast_2352_inst_req_1 : boolean;
  signal type_cast_2352_inst_ack_1 : boolean;
  signal phi_stmt_2349_req_0 : boolean;
  signal type_cast_2359_inst_req_0 : boolean;
  signal type_cast_2359_inst_ack_0 : boolean;
  signal type_cast_2359_inst_req_1 : boolean;
  signal type_cast_2359_inst_ack_1 : boolean;
  signal phi_stmt_2356_req_0 : boolean;
  signal phi_stmt_2335_ack_0 : boolean;
  signal phi_stmt_2342_ack_0 : boolean;
  signal phi_stmt_2349_ack_0 : boolean;
  signal phi_stmt_2356_ack_0 : boolean;
  signal phi_stmt_2543_req_1 : boolean;
  signal type_cast_2553_inst_req_0 : boolean;
  signal type_cast_2553_inst_ack_0 : boolean;
  signal type_cast_2553_inst_req_1 : boolean;
  signal type_cast_2553_inst_ack_1 : boolean;
  signal phi_stmt_2550_req_0 : boolean;
  signal type_cast_2559_inst_req_0 : boolean;
  signal type_cast_2559_inst_ack_0 : boolean;
  signal type_cast_2559_inst_req_1 : boolean;
  signal type_cast_2559_inst_ack_1 : boolean;
  signal phi_stmt_2556_req_0 : boolean;
  signal type_cast_2546_inst_req_0 : boolean;
  signal type_cast_2546_inst_ack_0 : boolean;
  signal type_cast_2546_inst_req_1 : boolean;
  signal type_cast_2546_inst_ack_1 : boolean;
  signal phi_stmt_2543_req_0 : boolean;
  signal type_cast_2555_inst_req_0 : boolean;
  signal type_cast_2555_inst_ack_0 : boolean;
  signal type_cast_2555_inst_req_1 : boolean;
  signal type_cast_2555_inst_ack_1 : boolean;
  signal phi_stmt_2550_req_1 : boolean;
  signal type_cast_2561_inst_req_0 : boolean;
  signal type_cast_2561_inst_ack_0 : boolean;
  signal type_cast_2561_inst_req_1 : boolean;
  signal type_cast_2561_inst_ack_1 : boolean;
  signal phi_stmt_2556_req_1 : boolean;
  signal phi_stmt_2543_ack_0 : boolean;
  signal phi_stmt_2550_ack_0 : boolean;
  signal phi_stmt_2556_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5768_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5768_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5768_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5768_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5768: Block -- control-path 
    signal convTransposeC_CP_5768_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5768_elements(0) <= convTransposeC_CP_5768_start;
    convTransposeC_CP_5768_symbol <= convTransposeC_CP_5768_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2209/$entry
      -- CP-element group 0: 	 branch_block_stmt_2209/branch_block_stmt_2209__entry__
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270__entry__
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/$entry
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_Sample/rr
      -- 
    cr_5961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(0), ack => type_cast_2242_inst_req_1); -- 
    cr_5989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(0), ack => type_cast_2255_inst_req_1); -- 
    rr_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(0), ack => RPIPE_Block2_start_2211_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2209/merge_stmt_2542__exit__
      -- CP-element group 1: 	 branch_block_stmt_2209/assign_stmt_2568__entry__
      -- CP-element group 1: 	 branch_block_stmt_2209/assign_stmt_2568__exit__
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2209/assign_stmt_2568/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/assign_stmt_2568/$exit
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/Update/cr
      -- 
    rr_6517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2341_inst_req_0); -- 
    cr_6522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2341_inst_req_1); -- 
    rr_6540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2348_inst_req_0); -- 
    cr_6545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2348_inst_req_1); -- 
    rr_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2352_inst_req_0); -- 
    cr_6568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2352_inst_req_1); -- 
    rr_6586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2359_inst_req_0); -- 
    cr_6591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(1), ack => type_cast_2359_inst_req_1); -- 
    convTransposeC_CP_5768_elements(1) <= convTransposeC_CP_5768_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_Update/cr
      -- 
    ra_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2211_inst_ack_0, ack => convTransposeC_CP_5768_elements(2)); -- 
    cr_5821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(2), ack => RPIPE_Block2_start_2211_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2211_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_Sample/rr
      -- 
    ca_5822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2211_inst_ack_1, ack => convTransposeC_CP_5768_elements(3)); -- 
    rr_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(3), ack => RPIPE_Block2_start_2214_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_Update/cr
      -- 
    ra_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2214_inst_ack_0, ack => convTransposeC_CP_5768_elements(4)); -- 
    cr_5835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(4), ack => RPIPE_Block2_start_2214_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2214_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_Sample/rr
      -- 
    ca_5836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2214_inst_ack_1, ack => convTransposeC_CP_5768_elements(5)); -- 
    rr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(5), ack => RPIPE_Block2_start_2217_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_Update/cr
      -- 
    ra_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2217_inst_ack_0, ack => convTransposeC_CP_5768_elements(6)); -- 
    cr_5849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(6), ack => RPIPE_Block2_start_2217_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2217_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_Sample/rr
      -- 
    ca_5850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2217_inst_ack_1, ack => convTransposeC_CP_5768_elements(7)); -- 
    rr_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(7), ack => RPIPE_Block2_start_2220_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_Update/$entry
      -- 
    ra_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2220_inst_ack_0, ack => convTransposeC_CP_5768_elements(8)); -- 
    cr_5863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(8), ack => RPIPE_Block2_start_2220_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2220_Update/$exit
      -- 
    ca_5864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2220_inst_ack_1, ack => convTransposeC_CP_5768_elements(9)); -- 
    rr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(9), ack => RPIPE_Block2_start_2223_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_Update/cr
      -- 
    ra_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2223_inst_ack_0, ack => convTransposeC_CP_5768_elements(10)); -- 
    cr_5877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(10), ack => RPIPE_Block2_start_2223_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2223_Update/ca
      -- 
    ca_5878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2223_inst_ack_1, ack => convTransposeC_CP_5768_elements(11)); -- 
    rr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(11), ack => RPIPE_Block2_start_2226_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_sample_completed_
      -- 
    ra_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2226_inst_ack_0, ack => convTransposeC_CP_5768_elements(12)); -- 
    cr_5891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(12), ack => RPIPE_Block2_start_2226_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2226_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_sample_start_
      -- 
    ca_5892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2226_inst_ack_1, ack => convTransposeC_CP_5768_elements(13)); -- 
    rr_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(13), ack => RPIPE_Block2_start_2229_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_Sample/ra
      -- 
    ra_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2229_inst_ack_0, ack => convTransposeC_CP_5768_elements(14)); -- 
    cr_5905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(14), ack => RPIPE_Block2_start_2229_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2229_Update/ca
      -- 
    ca_5906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2229_inst_ack_1, ack => convTransposeC_CP_5768_elements(15)); -- 
    rr_5914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(15), ack => RPIPE_Block2_start_2232_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_Update/cr
      -- 
    ra_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2232_inst_ack_0, ack => convTransposeC_CP_5768_elements(16)); -- 
    cr_5919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(16), ack => RPIPE_Block2_start_2232_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2232_Update/ca
      -- 
    ca_5920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2232_inst_ack_1, ack => convTransposeC_CP_5768_elements(17)); -- 
    rr_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(17), ack => RPIPE_Block2_start_2235_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_Update/$entry
      -- 
    ra_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2235_inst_ack_0, ack => convTransposeC_CP_5768_elements(18)); -- 
    cr_5933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(18), ack => RPIPE_Block2_start_2235_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2235_Update/$exit
      -- 
    ca_5934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2235_inst_ack_1, ack => convTransposeC_CP_5768_elements(19)); -- 
    rr_5942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(19), ack => RPIPE_Block2_start_2238_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_sample_completed_
      -- 
    ra_5943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2238_inst_ack_0, ack => convTransposeC_CP_5768_elements(20)); -- 
    cr_5947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(20), ack => RPIPE_Block2_start_2238_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2238_Update/ca
      -- 
    ca_5948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2238_inst_ack_1, ack => convTransposeC_CP_5768_elements(21)); -- 
    rr_5956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(21), ack => type_cast_2242_inst_req_0); -- 
    rr_5970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(21), ack => RPIPE_Block2_start_2251_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_Sample/$exit
      -- 
    ra_5957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2242_inst_ack_0, ack => convTransposeC_CP_5768_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2242_Update/ca
      -- 
    ca_5962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2242_inst_ack_1, ack => convTransposeC_CP_5768_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_Update/cr
      -- 
    ra_5971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2251_inst_ack_0, ack => convTransposeC_CP_5768_elements(24)); -- 
    cr_5975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(24), ack => RPIPE_Block2_start_2251_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2251_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_Sample/$entry
      -- 
    ca_5976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2251_inst_ack_1, ack => convTransposeC_CP_5768_elements(25)); -- 
    rr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(25), ack => type_cast_2255_inst_req_0); -- 
    rr_5998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(25), ack => RPIPE_Block2_start_2263_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_Sample/$exit
      -- 
    ra_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2255_inst_ack_0, ack => convTransposeC_CP_5768_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/type_cast_2255_update_completed_
      -- 
    ca_5990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2255_inst_ack_1, ack => convTransposeC_CP_5768_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_update_start_
      -- 
    ra_5999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2263_inst_ack_0, ack => convTransposeC_CP_5768_elements(28)); -- 
    cr_6003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(28), ack => RPIPE_Block2_start_2263_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2263_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_Sample/$entry
      -- 
    ca_6004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2263_inst_ack_1, ack => convTransposeC_CP_5768_elements(29)); -- 
    rr_6012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(29), ack => RPIPE_Block2_start_2266_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_Update/cr
      -- 
    ra_6013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2266_inst_ack_0, ack => convTransposeC_CP_5768_elements(30)); -- 
    cr_6017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(30), ack => RPIPE_Block2_start_2266_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2266_update_completed_
      -- 
    ca_6018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2266_inst_ack_1, ack => convTransposeC_CP_5768_elements(31)); -- 
    rr_6026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(31), ack => RPIPE_Block2_start_2269_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_Update/cr
      -- 
    ra_6027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2269_inst_ack_0, ack => convTransposeC_CP_5768_elements(32)); -- 
    cr_6031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(32), ack => RPIPE_Block2_start_2269_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/RPIPE_Block2_start_2269_update_completed_
      -- 
    ca_6032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2269_inst_ack_1, ack => convTransposeC_CP_5768_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270__exit__
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332__entry__
      -- CP-element group 34: 	 branch_block_stmt_2209/assign_stmt_2212_to_assign_stmt_2270/$exit
      -- 
    rr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2310_inst_req_0); -- 
    cr_6048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2302_inst_req_1); -- 
    cr_6090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2314_inst_req_1); -- 
    rr_6085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2314_inst_req_0); -- 
    cr_6062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2306_inst_req_1); -- 
    rr_6043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2302_inst_req_0); -- 
    cr_6076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2310_inst_req_1); -- 
    rr_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(34), ack => type_cast_2306_inst_req_0); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(23) & convTransposeC_CP_5768_elements(27) & convTransposeC_CP_5768_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_Sample/$exit
      -- 
    ra_6044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2302_inst_ack_0, ack => convTransposeC_CP_5768_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2302_Update/$exit
      -- 
    ca_6049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2302_inst_ack_1, ack => convTransposeC_CP_5768_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_Sample/$exit
      -- 
    ra_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_0, ack => convTransposeC_CP_5768_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2306_Update/ca
      -- 
    ca_6063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_1, ack => convTransposeC_CP_5768_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_sample_completed_
      -- 
    ra_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2310_inst_ack_0, ack => convTransposeC_CP_5768_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2310_update_completed_
      -- 
    ca_6077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2310_inst_ack_1, ack => convTransposeC_CP_5768_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_sample_completed_
      -- 
    ra_6086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2314_inst_ack_0, ack => convTransposeC_CP_5768_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/type_cast_2314_update_completed_
      -- 
    ca_6091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2314_inst_ack_1, ack => convTransposeC_CP_5768_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332/$exit
      -- CP-element group 43: 	 branch_block_stmt_2209/assign_stmt_2277_to_assign_stmt_2332__exit__
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2335/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2342/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2349/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/Update/cr
      -- 
    rr_6491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(43), ack => type_cast_2361_inst_req_0); -- 
    cr_6496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(43), ack => type_cast_2361_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(36) & convTransposeC_CP_5768_elements(38) & convTransposeC_CP_5768_elements(40) & convTransposeC_CP_5768_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_sample_completed_
      -- 
    ra_6103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2396_inst_ack_0, ack => convTransposeC_CP_5768_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_Update/ca
      -- 
    ca_6108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2396_inst_ack_1, ack => convTransposeC_CP_5768_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_Sample/ra
      -- 
    ra_6117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2400_inst_ack_0, ack => convTransposeC_CP_5768_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_Update/ca
      -- 
    ca_6122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2400_inst_ack_1, ack => convTransposeC_CP_5768_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_Sample/ra
      -- 
    ra_6131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_0, ack => convTransposeC_CP_5768_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_Update/ca
      -- 
    ca_6136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_1, ack => convTransposeC_CP_5768_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_Sample/ra
      -- 
    ra_6145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2434_inst_ack_0, ack => convTransposeC_CP_5768_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_Sample/req
      -- 
    ca_6150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2434_inst_ack_1, ack => convTransposeC_CP_5768_elements(51)); -- 
    req_6175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(51), ack => array_obj_ref_2440_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_Sample/ack
      -- 
    ack_6176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2440_index_offset_ack_0, ack => convTransposeC_CP_5768_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_request/req
      -- 
    ack_6181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2440_index_offset_ack_1, ack => convTransposeC_CP_5768_elements(53)); -- 
    req_6190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(53), ack => addr_of_2441_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_request/ack
      -- 
    ack_6191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2441_final_reg_ack_0, ack => convTransposeC_CP_5768_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Sample/word_access_start/word_0/rr
      -- 
    ack_6196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2441_final_reg_ack_1, ack => convTransposeC_CP_5768_elements(55)); -- 
    rr_6229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(55), ack => ptr_deref_2445_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Sample/word_access_start/word_0/ra
      -- 
    ra_6230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2445_load_0_ack_0, ack => convTransposeC_CP_5768_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/ptr_deref_2445_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/ptr_deref_2445_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/ptr_deref_2445_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/ptr_deref_2445_Merge/merge_ack
      -- 
    ca_6241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2445_load_0_ack_1, ack => convTransposeC_CP_5768_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_Sample/req
      -- 
    req_6271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(58), ack => array_obj_ref_2463_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(45) & convTransposeC_CP_5768_elements(47) & convTransposeC_CP_5768_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_Sample/ack
      -- 
    ack_6272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2463_index_offset_ack_0, ack => convTransposeC_CP_5768_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_request/req
      -- 
    ack_6277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2463_index_offset_ack_1, ack => convTransposeC_CP_5768_elements(60)); -- 
    req_6286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(60), ack => addr_of_2464_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_request/ack
      -- 
    ack_6287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2464_final_reg_ack_0, ack => convTransposeC_CP_5768_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_word_addrgen/root_register_ack
      -- 
    ack_6292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2464_final_reg_ack_1, ack => convTransposeC_CP_5768_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/ptr_deref_2467_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/ptr_deref_2467_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/ptr_deref_2467_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/ptr_deref_2467_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/word_access_start/word_0/rr
      -- 
    rr_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(63), ack => ptr_deref_2467_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(57) & convTransposeC_CP_5768_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Sample/word_access_start/word_0/ra
      -- 
    ra_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_store_0_ack_0, ack => convTransposeC_CP_5768_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Update/word_access_complete/word_0/ca
      -- 
    ca_6342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_store_0_ack_1, ack => convTransposeC_CP_5768_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_Sample/ra
      -- 
    ra_6351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2472_inst_ack_0, ack => convTransposeC_CP_5768_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_Update/ca
      -- 
    ca_6356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2472_inst_ack_1, ack => convTransposeC_CP_5768_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/$exit
      -- CP-element group 68: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484__exit__
      -- CP-element group 68: 	 branch_block_stmt_2209/if_stmt_2485__entry__
      -- CP-element group 68: 	 branch_block_stmt_2209/if_stmt_2485_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2209/if_stmt_2485_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2209/if_stmt_2485_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2209/if_stmt_2485_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2209/R_cmp_2486_place
      -- CP-element group 68: 	 branch_block_stmt_2209/if_stmt_2485_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2209/if_stmt_2485_else_link/$entry
      -- 
    branch_req_6364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(68), ack => if_stmt_2485_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(52) & convTransposeC_CP_5768_elements(59) & convTransposeC_CP_5768_elements(65) & convTransposeC_CP_5768_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2209/merge_stmt_2491__exit__
      -- CP-element group 69: 	 branch_block_stmt_2209/assign_stmt_2497__entry__
      -- CP-element group 69: 	 branch_block_stmt_2209/assign_stmt_2497__exit__
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2209/if_stmt_2485_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2209/if_stmt_2485_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2209/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2209/assign_stmt_2497/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/assign_stmt_2497/$exit
      -- CP-element group 69: 	 branch_block_stmt_2209/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2209/merge_stmt_2491_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2209/merge_stmt_2491_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/merge_stmt_2491_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2209/merge_stmt_2491_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2485_branch_ack_1, ack => convTransposeC_CP_5768_elements(69)); -- 
    rr_6701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2546_inst_req_0); -- 
    cr_6706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2546_inst_req_1); -- 
    rr_6724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2555_inst_req_0); -- 
    cr_6729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2555_inst_req_1); -- 
    rr_6747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2561_inst_req_0); -- 
    cr_6752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(69), ack => type_cast_2561_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2209/merge_stmt_2499__exit__
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535__entry__
      -- CP-element group 70: 	 branch_block_stmt_2209/if_stmt_2485_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2209/if_stmt_2485_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2209/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/$entry
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2209/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2209/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2209/merge_stmt_2499_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2209/merge_stmt_2499_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2209/merge_stmt_2499_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2209/merge_stmt_2499_PhiAck/dummy
      -- 
    else_choice_transition_6373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2485_branch_ack_0, ack => convTransposeC_CP_5768_elements(70)); -- 
    rr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(70), ack => type_cast_2513_inst_req_0); -- 
    cr_6394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(70), ack => type_cast_2513_inst_req_1); -- 
    cr_6408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(70), ack => type_cast_2529_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_Sample/ra
      -- 
    ra_6390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2513_inst_ack_0, ack => convTransposeC_CP_5768_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2513_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_Sample/rr
      -- 
    ca_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2513_inst_ack_1, ack => convTransposeC_CP_5768_elements(72)); -- 
    rr_6403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(72), ack => type_cast_2529_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_Sample/ra
      -- 
    ra_6404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2529_inst_ack_0, ack => convTransposeC_CP_5768_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535__exit__
      -- CP-element group 74: 	 branch_block_stmt_2209/if_stmt_2536__entry__
      -- CP-element group 74: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/$exit
      -- CP-element group 74: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2209/assign_stmt_2505_to_assign_stmt_2535/type_cast_2529_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2209/if_stmt_2536_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2209/if_stmt_2536_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2209/if_stmt_2536_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2209/if_stmt_2536_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2209/R_cmp122_2537_place
      -- CP-element group 74: 	 branch_block_stmt_2209/if_stmt_2536_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2209/if_stmt_2536_else_link/$entry
      -- 
    ca_6409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2529_inst_ack_1, ack => convTransposeC_CP_5768_elements(74)); -- 
    branch_req_6417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(74), ack => if_stmt_2536_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2209/merge_stmt_2570__exit__
      -- CP-element group 75: 	 branch_block_stmt_2209/assign_stmt_2575__entry__
      -- CP-element group 75: 	 branch_block_stmt_2209/if_stmt_2536_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2209/if_stmt_2536_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2209/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2209/assign_stmt_2575/$entry
      -- CP-element group 75: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2209/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2209/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2209/merge_stmt_2570_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2209/merge_stmt_2570_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2209/merge_stmt_2570_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2209/merge_stmt_2570_PhiAck/dummy
      -- 
    if_choice_transition_6422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2536_branch_ack_1, ack => convTransposeC_CP_5768_elements(75)); -- 
    req_6442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(75), ack => WPIPE_Block2_done_2572_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2209/if_stmt_2536_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2209/if_stmt_2536_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2543/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2536_branch_ack_0, ack => convTransposeC_CP_5768_elements(76)); -- 
    rr_6652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(76), ack => type_cast_2553_inst_req_0); -- 
    cr_6657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(76), ack => type_cast_2553_inst_req_1); -- 
    rr_6675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(76), ack => type_cast_2559_inst_req_0); -- 
    cr_6680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(76), ack => type_cast_2559_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_Update/req
      -- 
    ack_6443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2572_inst_ack_0, ack => convTransposeC_CP_5768_elements(77)); -- 
    req_6447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(77), ack => WPIPE_Block2_done_2572_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2209/$exit
      -- CP-element group 78: 	 branch_block_stmt_2209/branch_block_stmt_2209__exit__
      -- CP-element group 78: 	 branch_block_stmt_2209/assign_stmt_2575__exit__
      -- CP-element group 78: 	 branch_block_stmt_2209/return__
      -- CP-element group 78: 	 branch_block_stmt_2209/merge_stmt_2577__exit__
      -- CP-element group 78: 	 branch_block_stmt_2209/assign_stmt_2575/$exit
      -- CP-element group 78: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2209/assign_stmt_2575/WPIPE_Block2_done_2572_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2209/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2209/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2209/merge_stmt_2577_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2209/merge_stmt_2577_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2209/merge_stmt_2577_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2209/merge_stmt_2577_PhiAck/dummy
      -- 
    ack_6448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2572_inst_ack_1, ack => convTransposeC_CP_5768_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2335/$exit
      -- CP-element group 79: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2339_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_req
      -- 
    phi_stmt_2335_req_6459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2335_req_6459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(79), ack => phi_stmt_2335_req_0); -- 
    -- Element group convTransposeC_CP_5768_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5768_elements(43), ack => convTransposeC_CP_5768_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2342/$exit
      -- CP-element group 80: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2346_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_req
      -- 
    phi_stmt_2342_req_6467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2342_req_6467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(80), ack => phi_stmt_2342_req_0); -- 
    -- Element group convTransposeC_CP_5768_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5768_elements(43), ack => convTransposeC_CP_5768_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2349/$exit
      -- CP-element group 81: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2355_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_req
      -- 
    phi_stmt_2349_req_6475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2349_req_6475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(81), ack => phi_stmt_2349_req_1); -- 
    -- Element group convTransposeC_CP_5768_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeC_CP_5768_elements(43), ack => convTransposeC_CP_5768_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/Sample/ra
      -- 
    ra_6492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2361_inst_ack_0, ack => convTransposeC_CP_5768_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/Update/ca
      -- 
    ca_6497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2361_inst_ack_1, ack => convTransposeC_CP_5768_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/$exit
      -- CP-element group 84: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/$exit
      -- CP-element group 84: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2361/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_req
      -- 
    phi_stmt_2356_req_6498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2356_req_6498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(84), ack => phi_stmt_2356_req_1); -- 
    convTransposeC_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(82) & convTransposeC_CP_5768_elements(83);
      gj_convTransposeC_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2209/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(79) & convTransposeC_CP_5768_elements(80) & convTransposeC_CP_5768_elements(81) & convTransposeC_CP_5768_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/Sample/ra
      -- 
    ra_6518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_0, ack => convTransposeC_CP_5768_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/Update/ca
      -- 
    ca_6523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_1, ack => convTransposeC_CP_5768_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/$exit
      -- CP-element group 88: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/$exit
      -- CP-element group 88: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_sources/type_cast_2341/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2335/phi_stmt_2335_req
      -- 
    phi_stmt_2335_req_6524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2335_req_6524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(88), ack => phi_stmt_2335_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(86) & convTransposeC_CP_5768_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/Sample/ra
      -- 
    ra_6541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2348_inst_ack_0, ack => convTransposeC_CP_5768_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/Update/ca
      -- 
    ca_6546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2348_inst_ack_1, ack => convTransposeC_CP_5768_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/$exit
      -- CP-element group 91: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/$exit
      -- CP-element group 91: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_sources/type_cast_2348/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2342/phi_stmt_2342_req
      -- 
    phi_stmt_2342_req_6547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2342_req_6547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(91), ack => phi_stmt_2342_req_1); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(89) & convTransposeC_CP_5768_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/Sample/ra
      -- 
    ra_6564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_0, ack => convTransposeC_CP_5768_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/Update/ca
      -- 
    ca_6569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_1, ack => convTransposeC_CP_5768_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/$exit
      -- CP-element group 94: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/$exit
      -- CP-element group 94: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_sources/type_cast_2352/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2349/phi_stmt_2349_req
      -- 
    phi_stmt_2349_req_6570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2349_req_6570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(94), ack => phi_stmt_2349_req_0); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(92) & convTransposeC_CP_5768_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/Sample/ra
      -- 
    ra_6587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2359_inst_ack_0, ack => convTransposeC_CP_5768_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/Update/ca
      -- 
    ca_6592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2359_inst_ack_1, ack => convTransposeC_CP_5768_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/$exit
      -- CP-element group 97: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/$exit
      -- CP-element group 97: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_sources/type_cast_2359/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2356/phi_stmt_2356_req
      -- 
    phi_stmt_2356_req_6593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2356_req_6593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(97), ack => phi_stmt_2356_req_0); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(95) & convTransposeC_CP_5768_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2209/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(88) & convTransposeC_CP_5768_elements(91) & convTransposeC_CP_5768_elements(94) & convTransposeC_CP_5768_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2209/merge_stmt_2334_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2209/merge_stmt_2334_PhiAck/$entry
      -- 
    convTransposeC_CP_5768_elements(99) <= OrReduce(convTransposeC_CP_5768_elements(85) & convTransposeC_CP_5768_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2209/merge_stmt_2334_PhiAck/phi_stmt_2335_ack
      -- 
    phi_stmt_2335_ack_6598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2335_ack_0, ack => convTransposeC_CP_5768_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2209/merge_stmt_2334_PhiAck/phi_stmt_2342_ack
      -- 
    phi_stmt_2342_ack_6599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2342_ack_0, ack => convTransposeC_CP_5768_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2209/merge_stmt_2334_PhiAck/phi_stmt_2349_ack
      -- 
    phi_stmt_2349_ack_6600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2349_ack_0, ack => convTransposeC_CP_5768_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2209/merge_stmt_2334_PhiAck/phi_stmt_2356_ack
      -- 
    phi_stmt_2356_ack_6601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2356_ack_0, ack => convTransposeC_CP_5768_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2396_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2209/merge_stmt_2334__exit__
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484__entry__
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2400_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2404_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2434_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2440_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2441_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2445_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/array_obj_ref_2463_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/addr_of_2464_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/ptr_deref_2467_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2209/assign_stmt_2368_to_assign_stmt_2484/type_cast_2472_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2209/merge_stmt_2334_PhiAck/$exit
      -- 
    rr_6102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2396_inst_req_0); -- 
    cr_6107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2396_inst_req_1); -- 
    rr_6116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2400_inst_req_0); -- 
    cr_6121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2400_inst_req_1); -- 
    rr_6130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2404_inst_req_0); -- 
    cr_6135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2404_inst_req_1); -- 
    rr_6144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2434_inst_req_0); -- 
    cr_6149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2434_inst_req_1); -- 
    req_6180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => array_obj_ref_2440_index_offset_req_1); -- 
    req_6195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => addr_of_2441_final_reg_req_1); -- 
    cr_6240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => ptr_deref_2445_load_0_req_1); -- 
    req_6276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => array_obj_ref_2463_index_offset_req_1); -- 
    req_6291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => addr_of_2464_final_reg_req_1); -- 
    cr_6341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => ptr_deref_2467_store_0_req_1); -- 
    rr_6350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2472_inst_req_0); -- 
    cr_6355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(104), ack => type_cast_2472_inst_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(100) & convTransposeC_CP_5768_elements(101) & convTransposeC_CP_5768_elements(102) & convTransposeC_CP_5768_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2543/$exit
      -- CP-element group 105: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2549_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_req
      -- 
    phi_stmt_2543_req_6636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2543_req_6636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(105), ack => phi_stmt_2543_req_1); -- 
    -- Element group convTransposeC_CP_5768_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5768_elements(76), ack => convTransposeC_CP_5768_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/Sample/ra
      -- 
    ra_6653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2553_inst_ack_0, ack => convTransposeC_CP_5768_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/Update/ca
      -- 
    ca_6658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2553_inst_ack_1, ack => convTransposeC_CP_5768_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/$exit
      -- CP-element group 108: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/$exit
      -- CP-element group 108: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2553/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_req
      -- 
    phi_stmt_2550_req_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2550_req_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(108), ack => phi_stmt_2550_req_0); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(106) & convTransposeC_CP_5768_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Sample/ra
      -- 
    ra_6676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_0, ack => convTransposeC_CP_5768_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/Update/ca
      -- 
    ca_6681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_1, ack => convTransposeC_CP_5768_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/$exit
      -- CP-element group 111: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/$exit
      -- CP-element group 111: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2559/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_req
      -- 
    phi_stmt_2556_req_6682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2556_req_6682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(111), ack => phi_stmt_2556_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(109) & convTransposeC_CP_5768_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2209/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(105) & convTransposeC_CP_5768_elements(108) & convTransposeC_CP_5768_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Sample/ra
      -- 
    ra_6702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2546_inst_ack_0, ack => convTransposeC_CP_5768_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/Update/ca
      -- 
    ca_6707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2546_inst_ack_1, ack => convTransposeC_CP_5768_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/$exit
      -- CP-element group 115: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/$exit
      -- CP-element group 115: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_sources/type_cast_2546/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2543/phi_stmt_2543_req
      -- 
    phi_stmt_2543_req_6708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2543_req_6708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(115), ack => phi_stmt_2543_req_0); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(113) & convTransposeC_CP_5768_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/Sample/ra
      -- 
    ra_6725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2555_inst_ack_0, ack => convTransposeC_CP_5768_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/Update/ca
      -- 
    ca_6730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2555_inst_ack_1, ack => convTransposeC_CP_5768_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/$exit
      -- CP-element group 118: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/$exit
      -- CP-element group 118: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_sources/type_cast_2555/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2550/phi_stmt_2550_req
      -- 
    phi_stmt_2550_req_6731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2550_req_6731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(118), ack => phi_stmt_2550_req_1); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(116) & convTransposeC_CP_5768_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Sample/ra
      -- 
    ra_6748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2561_inst_ack_0, ack => convTransposeC_CP_5768_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/Update/ca
      -- 
    ca_6753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2561_inst_ack_1, ack => convTransposeC_CP_5768_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/$exit
      -- CP-element group 121: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/$exit
      -- CP-element group 121: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_sources/type_cast_2561/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2556/phi_stmt_2556_req
      -- 
    phi_stmt_2556_req_6754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2556_req_6754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5768_elements(121), ack => phi_stmt_2556_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(119) & convTransposeC_CP_5768_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2209/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(115) & convTransposeC_CP_5768_elements(118) & convTransposeC_CP_5768_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2209/merge_stmt_2542_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2209/merge_stmt_2542_PhiAck/$entry
      -- 
    convTransposeC_CP_5768_elements(123) <= OrReduce(convTransposeC_CP_5768_elements(112) & convTransposeC_CP_5768_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2209/merge_stmt_2542_PhiAck/phi_stmt_2543_ack
      -- 
    phi_stmt_2543_ack_6759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2543_ack_0, ack => convTransposeC_CP_5768_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2209/merge_stmt_2542_PhiAck/phi_stmt_2550_ack
      -- 
    phi_stmt_2550_ack_6760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2550_ack_0, ack => convTransposeC_CP_5768_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2209/merge_stmt_2542_PhiAck/phi_stmt_2556_ack
      -- 
    phi_stmt_2556_ack_6761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2556_ack_0, ack => convTransposeC_CP_5768_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2209/merge_stmt_2542_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5768_elements(124) & convTransposeC_CP_5768_elements(125) & convTransposeC_CP_5768_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5768_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2462_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2462_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2439_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2439_scaled : std_logic_vector(13 downto 0);
    signal add121_2332 : std_logic_vector(31 downto 0);
    signal add45_2283 : std_logic_vector(15 downto 0);
    signal add58_2294 : std_logic_vector(15 downto 0);
    signal add77_2415 : std_logic_vector(63 downto 0);
    signal add79_2425 : std_logic_vector(63 downto 0);
    signal add91_2479 : std_logic_vector(31 downto 0);
    signal add98_2497 : std_logic_vector(15 downto 0);
    signal add_2261 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2373 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2440_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2440_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2440_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2440_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2440_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2440_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2463_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2463_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2463_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2463_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2463_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2463_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2442 : std_logic_vector(31 downto 0);
    signal arrayidx87_2465 : std_logic_vector(31 downto 0);
    signal call11_2230 : std_logic_vector(15 downto 0);
    signal call13_2233 : std_logic_vector(15 downto 0);
    signal call14_2236 : std_logic_vector(15 downto 0);
    signal call15_2239 : std_logic_vector(15 downto 0);
    signal call16_2252 : std_logic_vector(15 downto 0);
    signal call18_2264 : std_logic_vector(15 downto 0);
    signal call1_2215 : std_logic_vector(15 downto 0);
    signal call20_2267 : std_logic_vector(15 downto 0);
    signal call22_2270 : std_logic_vector(15 downto 0);
    signal call3_2218 : std_logic_vector(15 downto 0);
    signal call5_2221 : std_logic_vector(15 downto 0);
    signal call7_2224 : std_logic_vector(15 downto 0);
    signal call9_2227 : std_logic_vector(15 downto 0);
    signal call_2212 : std_logic_vector(15 downto 0);
    signal cmp106_2510 : std_logic_vector(0 downto 0);
    signal cmp122_2535 : std_logic_vector(0 downto 0);
    signal cmp_2484 : std_logic_vector(0 downto 0);
    signal conv112_2530 : std_logic_vector(31 downto 0);
    signal conv115_2315 : std_logic_vector(31 downto 0);
    signal conv17_2256 : std_logic_vector(31 downto 0);
    signal conv65_2397 : std_logic_vector(63 downto 0);
    signal conv68_2303 : std_logic_vector(63 downto 0);
    signal conv70_2401 : std_logic_vector(63 downto 0);
    signal conv73_2307 : std_logic_vector(63 downto 0);
    signal conv75_2405 : std_logic_vector(63 downto 0);
    signal conv90_2473 : std_logic_vector(31 downto 0);
    signal conv94_2311 : std_logic_vector(31 downto 0);
    signal conv_2243 : std_logic_vector(31 downto 0);
    signal idxprom86_2458 : std_logic_vector(63 downto 0);
    signal idxprom_2435 : std_logic_vector(63 downto 0);
    signal inc110_2514 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2519 : std_logic_vector(15 downto 0);
    signal inc_2505 : std_logic_vector(15 downto 0);
    signal indvar_2335 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2568 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2556 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2356 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2550 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2349 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2526 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2543 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2342 : std_logic_vector(15 downto 0);
    signal mul54_2388 : std_logic_vector(15 downto 0);
    signal mul76_2410 : std_logic_vector(63 downto 0);
    signal mul78_2420 : std_logic_vector(63 downto 0);
    signal mul_2378 : std_logic_vector(15 downto 0);
    signal ptr_deref_2445_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2445_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2445_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2445_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2445_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2467_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2467_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2467_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2467_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2467_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2467_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2249 : std_logic_vector(31 downto 0);
    signal shr116137_2321 : std_logic_vector(31 downto 0);
    signal shr120138_2327 : std_logic_vector(31 downto 0);
    signal shr136_2277 : std_logic_vector(15 downto 0);
    signal shr81_2431 : std_logic_vector(31 downto 0);
    signal shr85_2452 : std_logic_vector(63 downto 0);
    signal sub48_2383 : std_logic_vector(15 downto 0);
    signal sub61_2299 : std_logic_vector(15 downto 0);
    signal sub62_2393 : std_logic_vector(15 downto 0);
    signal sub_2288 : std_logic_vector(15 downto 0);
    signal tmp1_2368 : std_logic_vector(31 downto 0);
    signal tmp83_2446 : std_logic_vector(63 downto 0);
    signal type_cast_2247_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2275_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2281_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2292_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2319_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2325_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2339_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2341_wire : std_logic_vector(31 downto 0);
    signal type_cast_2346_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2348_wire : std_logic_vector(15 downto 0);
    signal type_cast_2352_wire : std_logic_vector(15 downto 0);
    signal type_cast_2355_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2359_wire : std_logic_vector(15 downto 0);
    signal type_cast_2361_wire : std_logic_vector(15 downto 0);
    signal type_cast_2366_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2429_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2450_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2456_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2477_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2495_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2503_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2523_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2546_wire : std_logic_vector(15 downto 0);
    signal type_cast_2549_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2553_wire : std_logic_vector(15 downto 0);
    signal type_cast_2555_wire : std_logic_vector(15 downto 0);
    signal type_cast_2559_wire : std_logic_vector(15 downto 0);
    signal type_cast_2561_wire : std_logic_vector(15 downto 0);
    signal type_cast_2566_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2574_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2440_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2440_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2440_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2440_resized_base_address <= "00000000000000";
    array_obj_ref_2463_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2463_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2463_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2463_resized_base_address <= "00000000000000";
    ptr_deref_2445_word_offset_0 <= "00000000000000";
    ptr_deref_2467_word_offset_0 <= "00000000000000";
    type_cast_2247_wire_constant <= "00000000000000000000000000010000";
    type_cast_2275_wire_constant <= "0000000000000001";
    type_cast_2281_wire_constant <= "1111111111111111";
    type_cast_2292_wire_constant <= "1111111111111111";
    type_cast_2319_wire_constant <= "00000000000000000000000000000010";
    type_cast_2325_wire_constant <= "00000000000000000000000000000001";
    type_cast_2339_wire_constant <= "00000000000000000000000000000000";
    type_cast_2346_wire_constant <= "0000000000000000";
    type_cast_2355_wire_constant <= "0000000000000000";
    type_cast_2366_wire_constant <= "00000000000000000000000000000100";
    type_cast_2429_wire_constant <= "00000000000000000000000000000010";
    type_cast_2450_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2456_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2477_wire_constant <= "00000000000000000000000000000100";
    type_cast_2495_wire_constant <= "0000000000000100";
    type_cast_2503_wire_constant <= "0000000000000001";
    type_cast_2523_wire_constant <= "0000000000000000";
    type_cast_2549_wire_constant <= "0000000000000000";
    type_cast_2566_wire_constant <= "00000000000000000000000000000001";
    type_cast_2574_wire_constant <= "0000000000000001";
    phi_stmt_2335: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2339_wire_constant & type_cast_2341_wire;
      req <= phi_stmt_2335_req_0 & phi_stmt_2335_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2335",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2335_ack_0,
          idata => idata,
          odata => indvar_2335,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2335
    phi_stmt_2342: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2346_wire_constant & type_cast_2348_wire;
      req <= phi_stmt_2342_req_0 & phi_stmt_2342_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2342",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2342_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2342,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2342
    phi_stmt_2349: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2352_wire & type_cast_2355_wire_constant;
      req <= phi_stmt_2349_req_0 & phi_stmt_2349_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2349",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2349_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2349,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2349
    phi_stmt_2356: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2359_wire & type_cast_2361_wire;
      req <= phi_stmt_2356_req_0 & phi_stmt_2356_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2356",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2356_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2356,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2356
    phi_stmt_2543: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2546_wire & type_cast_2549_wire_constant;
      req <= phi_stmt_2543_req_0 & phi_stmt_2543_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2543",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2543_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2543,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2543
    phi_stmt_2550: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2553_wire & type_cast_2555_wire;
      req <= phi_stmt_2550_req_0 & phi_stmt_2550_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2550",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2550_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2550,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2550
    phi_stmt_2556: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2559_wire & type_cast_2561_wire;
      req <= phi_stmt_2556_req_0 & phi_stmt_2556_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2556",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2556_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2556,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2556
    -- flow-through select operator MUX_2525_inst
    input_dim1x_x2_2526 <= type_cast_2523_wire_constant when (cmp106_2510(0) /=  '0') else inc_2505;
    addr_of_2441_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2441_final_reg_req_0;
      addr_of_2441_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2441_final_reg_req_1;
      addr_of_2441_final_reg_ack_1<= rack(0);
      addr_of_2441_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2441_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2440_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2464_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2464_final_reg_req_0;
      addr_of_2464_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2464_final_reg_req_1;
      addr_of_2464_final_reg_ack_1<= rack(0);
      addr_of_2464_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2464_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2463_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2465,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2242_inst_req_0;
      type_cast_2242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2242_inst_req_1;
      type_cast_2242_inst_ack_1<= rack(0);
      type_cast_2242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2242_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2239,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2255_inst_req_0;
      type_cast_2255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2255_inst_req_1;
      type_cast_2255_inst_ack_1<= rack(0);
      type_cast_2255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2302_inst_req_0;
      type_cast_2302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2302_inst_req_1;
      type_cast_2302_inst_ack_1<= rack(0);
      type_cast_2302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2270,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2306_inst_req_0;
      type_cast_2306_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2306_inst_req_1;
      type_cast_2306_inst_ack_1<= rack(0);
      type_cast_2306_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2267,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2307,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2310_inst_req_0;
      type_cast_2310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2310_inst_req_1;
      type_cast_2310_inst_ack_1<= rack(0);
      type_cast_2310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2218,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2314_inst_req_0;
      type_cast_2314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2314_inst_req_1;
      type_cast_2314_inst_ack_1<= rack(0);
      type_cast_2314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2212,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2341_inst_req_0;
      type_cast_2341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2341_inst_req_1;
      type_cast_2341_inst_ack_1<= rack(0);
      type_cast_2341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2568,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2341_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2348_inst_req_0;
      type_cast_2348_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2348_inst_req_1;
      type_cast_2348_inst_ack_1<= rack(0);
      type_cast_2348_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2543,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2348_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2352_inst_req_0;
      type_cast_2352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2352_inst_req_1;
      type_cast_2352_inst_ack_1<= rack(0);
      type_cast_2352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2550,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2352_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2359_inst_req_0;
      type_cast_2359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2359_inst_req_1;
      type_cast_2359_inst_ack_1<= rack(0);
      type_cast_2359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2359_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2361_inst_req_0;
      type_cast_2361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2361_inst_req_1;
      type_cast_2361_inst_ack_1<= rack(0);
      type_cast_2361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2277,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2361_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2396_inst_req_0;
      type_cast_2396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2396_inst_req_1;
      type_cast_2396_inst_ack_1<= rack(0);
      type_cast_2396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2400_inst_req_0;
      type_cast_2400_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2400_inst_req_1;
      type_cast_2400_inst_ack_1<= rack(0);
      type_cast_2400_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2400_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2401,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2404_inst_req_0;
      type_cast_2404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2404_inst_req_1;
      type_cast_2404_inst_ack_1<= rack(0);
      type_cast_2404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2404_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2405,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2434_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2434_inst_req_0;
      type_cast_2434_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2434_inst_req_1;
      type_cast_2434_inst_ack_1<= rack(0);
      type_cast_2434_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2434_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2431,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2435,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2472_inst_req_0;
      type_cast_2472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2472_inst_req_1;
      type_cast_2472_inst_ack_1<= rack(0);
      type_cast_2472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2513_inst_req_0;
      type_cast_2513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2513_inst_req_1;
      type_cast_2513_inst_ack_1<= rack(0);
      type_cast_2513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2510,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2529_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2529_inst_req_0;
      type_cast_2529_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2529_inst_req_1;
      type_cast_2529_inst_ack_1<= rack(0);
      type_cast_2529_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2529_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2519,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2530,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2546_inst_req_0;
      type_cast_2546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2546_inst_req_1;
      type_cast_2546_inst_ack_1<= rack(0);
      type_cast_2546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2546_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2546_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2553_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2553_inst_req_0;
      type_cast_2553_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2553_inst_req_1;
      type_cast_2553_inst_ack_1<= rack(0);
      type_cast_2553_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2553_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2526,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2553_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2555_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2555_inst_req_0;
      type_cast_2555_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2555_inst_req_1;
      type_cast_2555_inst_ack_1<= rack(0);
      type_cast_2555_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2555_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2555_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2559_inst_req_0;
      type_cast_2559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2559_inst_req_1;
      type_cast_2559_inst_ack_1<= rack(0);
      type_cast_2559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2519,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2559_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2561_inst_req_0;
      type_cast_2561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2561_inst_req_1;
      type_cast_2561_inst_ack_1<= rack(0);
      type_cast_2561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2561_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2440_index_1_rename
    process(R_idxprom_2439_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2439_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2439_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2440_index_1_resize
    process(idxprom_2435) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2435;
      ov := iv(13 downto 0);
      R_idxprom_2439_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2440_root_address_inst
    process(array_obj_ref_2440_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2440_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2440_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2463_index_1_rename
    process(R_idxprom86_2462_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2462_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2462_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2463_index_1_resize
    process(idxprom86_2458) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2458;
      ov := iv(13 downto 0);
      R_idxprom86_2462_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2463_root_address_inst
    process(array_obj_ref_2463_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2463_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2463_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2445_addr_0
    process(ptr_deref_2445_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2445_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2445_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2445_base_resize
    process(arrayidx82_2442) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2442;
      ov := iv(13 downto 0);
      ptr_deref_2445_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2445_gather_scatter
    process(ptr_deref_2445_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2445_data_0;
      ov(63 downto 0) := iv;
      tmp83_2446 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2445_root_address_inst
    process(ptr_deref_2445_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2445_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2445_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2467_addr_0
    process(ptr_deref_2467_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2467_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2467_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2467_base_resize
    process(arrayidx87_2465) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2465;
      ov := iv(13 downto 0);
      ptr_deref_2467_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2467_gather_scatter
    process(tmp83_2446) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2446;
      ov(63 downto 0) := iv;
      ptr_deref_2467_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2467_root_address_inst
    process(ptr_deref_2467_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2467_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2467_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2485_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2484;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2485_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2485_branch_req_0,
          ack0 => if_stmt_2485_branch_ack_0,
          ack1 => if_stmt_2485_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2536_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2535;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2536_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2536_branch_req_0,
          ack0 => if_stmt_2536_branch_ack_0,
          ack1 => if_stmt_2536_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2282_inst
    process(call7_2224) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2224, type_cast_2281_wire_constant, tmp_var);
      add45_2283 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2293_inst
    process(call9_2227) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2227, type_cast_2292_wire_constant, tmp_var);
      add58_2294 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2382_inst
    process(sub_2288, mul_2378) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2288, mul_2378, tmp_var);
      sub48_2383 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2392_inst
    process(sub61_2299, mul54_2388) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2299, mul54_2388, tmp_var);
      sub62_2393 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2496_inst
    process(input_dim2x_x1_2342) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2342, type_cast_2495_wire_constant, tmp_var);
      add98_2497 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2504_inst
    process(input_dim1x_x1_2349) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2349, type_cast_2503_wire_constant, tmp_var);
      inc_2505 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2518_inst
    process(inc110_2514, input_dim0x_x2_2356) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2514, input_dim0x_x2_2356, tmp_var);
      inc110x_xinput_dim0x_x2_2519 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2331_inst
    process(shr116137_2321, shr120138_2327) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2321, shr120138_2327, tmp_var);
      add121_2332 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2372_inst
    process(add_2261, tmp1_2368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2261, tmp1_2368, tmp_var);
      add_src_0x_x0_2373 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2478_inst
    process(conv90_2473) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2473, type_cast_2477_wire_constant, tmp_var);
      add91_2479 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2567_inst
    process(indvar_2335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2335, type_cast_2566_wire_constant, tmp_var);
      indvarx_xnext_2568 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2414_inst
    process(mul76_2410, conv70_2401) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2410, conv70_2401, tmp_var);
      add77_2415 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2424_inst
    process(mul78_2420, conv65_2397) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2420, conv65_2397, tmp_var);
      add79_2425 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2457_inst
    process(shr85_2452) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2452, type_cast_2456_wire_constant, tmp_var);
      idxprom86_2458 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2509_inst
    process(inc_2505, call1_2215) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2505, call1_2215, tmp_var);
      cmp106_2510 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2534_inst
    process(conv112_2530, add121_2332) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2530, add121_2332, tmp_var);
      cmp122_2535 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2276_inst
    process(call_2212) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2212, type_cast_2275_wire_constant, tmp_var);
      shr136_2277 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2320_inst
    process(conv115_2315) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2315, type_cast_2319_wire_constant, tmp_var);
      shr116137_2321 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2326_inst
    process(conv115_2315) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2315, type_cast_2325_wire_constant, tmp_var);
      shr120138_2327 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2430_inst
    process(add_src_0x_x0_2373) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2373, type_cast_2429_wire_constant, tmp_var);
      shr81_2431 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2451_inst
    process(add79_2425) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2425, type_cast_2450_wire_constant, tmp_var);
      shr85_2452 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2377_inst
    process(input_dim0x_x2_2356, call13_2233) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2356, call13_2233, tmp_var);
      mul_2378 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2387_inst
    process(input_dim1x_x1_2349, call13_2233) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2349, call13_2233, tmp_var);
      mul54_2388 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2367_inst
    process(indvar_2335) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2335, type_cast_2366_wire_constant, tmp_var);
      tmp1_2368 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2409_inst
    process(conv75_2405, conv73_2307) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2405, conv73_2307, tmp_var);
      mul76_2410 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2419_inst
    process(add77_2415, conv68_2303) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2415, conv68_2303, tmp_var);
      mul78_2420 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2260_inst
    process(shl_2249, conv17_2256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2249, conv17_2256, tmp_var);
      add_2261 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2248_inst
    process(conv_2243) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2243, type_cast_2247_wire_constant, tmp_var);
      shl_2249 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2287_inst
    process(add45_2283, call14_2236) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2283, call14_2236, tmp_var);
      sub_2288 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2298_inst
    process(add58_2294, call14_2236) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2294, call14_2236, tmp_var);
      sub61_2299 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2483_inst
    process(add91_2479, conv94_2311) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2479, conv94_2311, tmp_var);
      cmp_2484 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2440_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2439_scaled;
      array_obj_ref_2440_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2440_index_offset_req_0;
      array_obj_ref_2440_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2440_index_offset_req_1;
      array_obj_ref_2440_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2463_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2462_scaled;
      array_obj_ref_2463_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2463_index_offset_req_0;
      array_obj_ref_2463_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2463_index_offset_req_1;
      array_obj_ref_2463_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2445_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2445_load_0_req_0;
      ptr_deref_2445_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2445_load_0_req_1;
      ptr_deref_2445_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2445_word_address_0;
      ptr_deref_2445_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2467_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2467_store_0_req_0;
      ptr_deref_2467_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2467_store_0_req_1;
      ptr_deref_2467_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2467_word_address_0;
      data_in <= ptr_deref_2467_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2251_inst RPIPE_Block2_start_2263_inst RPIPE_Block2_start_2266_inst RPIPE_Block2_start_2269_inst RPIPE_Block2_start_2238_inst RPIPE_Block2_start_2235_inst RPIPE_Block2_start_2232_inst RPIPE_Block2_start_2229_inst RPIPE_Block2_start_2226_inst RPIPE_Block2_start_2223_inst RPIPE_Block2_start_2220_inst RPIPE_Block2_start_2217_inst RPIPE_Block2_start_2214_inst RPIPE_Block2_start_2211_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2251_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2263_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2266_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2269_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2238_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2235_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2232_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2229_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2226_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2223_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2220_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2217_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2214_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2211_inst_req_0;
      RPIPE_Block2_start_2251_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2263_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2266_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2269_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2238_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2235_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2232_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2229_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2226_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2223_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2220_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2217_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2214_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2211_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2251_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2263_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2266_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2269_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2238_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2235_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2232_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2229_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2226_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2223_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2220_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2217_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2214_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2211_inst_req_1;
      RPIPE_Block2_start_2251_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2263_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2266_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2269_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2238_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2235_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2232_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2229_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2226_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2223_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2220_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2217_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2214_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2211_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call16_2252 <= data_out(223 downto 208);
      call18_2264 <= data_out(207 downto 192);
      call20_2267 <= data_out(191 downto 176);
      call22_2270 <= data_out(175 downto 160);
      call15_2239 <= data_out(159 downto 144);
      call14_2236 <= data_out(143 downto 128);
      call13_2233 <= data_out(127 downto 112);
      call11_2230 <= data_out(111 downto 96);
      call9_2227 <= data_out(95 downto 80);
      call7_2224 <= data_out(79 downto 64);
      call5_2221 <= data_out(63 downto 48);
      call3_2218 <= data_out(47 downto 32);
      call1_2215 <= data_out(31 downto 16);
      call_2212 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2572_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2572_inst_req_0;
      WPIPE_Block2_done_2572_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2572_inst_req_1;
      WPIPE_Block2_done_2572_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2574_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6778_start: Boolean;
  signal convTransposeD_CP_6778_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2592_inst_ack_1 : boolean;
  signal type_cast_2614_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2583_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2589_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2610_inst_ack_1 : boolean;
  signal type_cast_2627_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2604_inst_req_1 : boolean;
  signal type_cast_2627_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2583_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2583_inst_req_0 : boolean;
  signal type_cast_2689_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2589_inst_req_0 : boolean;
  signal type_cast_2689_inst_req_1 : boolean;
  signal type_cast_2693_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2595_inst_ack_1 : boolean;
  signal type_cast_2689_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2595_inst_req_1 : boolean;
  signal type_cast_2614_inst_ack_0 : boolean;
  signal type_cast_2685_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2601_inst_ack_1 : boolean;
  signal type_cast_2758_inst_req_0 : boolean;
  signal type_cast_2758_inst_ack_0 : boolean;
  signal type_cast_2758_inst_req_1 : boolean;
  signal type_cast_2758_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2601_inst_req_0 : boolean;
  signal type_cast_2685_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2583_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2638_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2607_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2607_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2592_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2623_inst_req_1 : boolean;
  signal type_cast_2693_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2623_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2623_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2638_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2592_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2589_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2623_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2604_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2586_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2601_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2601_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2595_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2607_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2586_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2610_inst_req_1 : boolean;
  signal type_cast_2614_inst_req_1 : boolean;
  signal type_cast_2614_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2592_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2641_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2638_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2641_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2604_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2635_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2635_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2586_inst_ack_0 : boolean;
  signal type_cast_2689_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2589_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2638_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2595_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2641_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2604_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2635_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2635_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2641_inst_ack_1 : boolean;
  signal type_cast_2685_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2586_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2607_inst_ack_1 : boolean;
  signal type_cast_2762_inst_req_1 : boolean;
  signal type_cast_2762_inst_ack_1 : boolean;
  signal type_cast_2766_inst_req_0 : boolean;
  signal type_cast_2627_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2610_inst_ack_0 : boolean;
  signal type_cast_2796_inst_req_0 : boolean;
  signal type_cast_2796_inst_ack_0 : boolean;
  signal type_cast_2796_inst_ack_1 : boolean;
  signal type_cast_2627_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2610_inst_req_0 : boolean;
  signal type_cast_2796_inst_req_1 : boolean;
  signal addr_of_2803_final_reg_req_0 : boolean;
  signal addr_of_2803_final_reg_ack_0 : boolean;
  signal addr_of_2803_final_reg_req_1 : boolean;
  signal addr_of_2803_final_reg_ack_1 : boolean;
  signal array_obj_ref_2802_index_offset_ack_0 : boolean;
  signal array_obj_ref_2802_index_offset_req_1 : boolean;
  signal array_obj_ref_2802_index_offset_ack_1 : boolean;
  signal RPIPE_Block3_start_2598_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2598_inst_req_1 : boolean;
  signal type_cast_2766_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2598_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2598_inst_req_0 : boolean;
  signal type_cast_2693_inst_ack_0 : boolean;
  signal type_cast_2766_inst_req_1 : boolean;
  signal type_cast_2766_inst_ack_1 : boolean;
  signal array_obj_ref_2802_index_offset_req_0 : boolean;
  signal type_cast_2762_inst_req_0 : boolean;
  signal type_cast_2762_inst_ack_0 : boolean;
  signal type_cast_2693_inst_req_0 : boolean;
  signal type_cast_2685_inst_ack_0 : boolean;
  signal ptr_deref_2807_load_0_req_0 : boolean;
  signal ptr_deref_2807_load_0_ack_0 : boolean;
  signal ptr_deref_2807_load_0_req_1 : boolean;
  signal ptr_deref_2807_load_0_ack_1 : boolean;
  signal array_obj_ref_2825_index_offset_req_0 : boolean;
  signal array_obj_ref_2825_index_offset_ack_0 : boolean;
  signal array_obj_ref_2825_index_offset_req_1 : boolean;
  signal array_obj_ref_2825_index_offset_ack_1 : boolean;
  signal addr_of_2826_final_reg_req_0 : boolean;
  signal addr_of_2826_final_reg_ack_0 : boolean;
  signal addr_of_2826_final_reg_req_1 : boolean;
  signal addr_of_2826_final_reg_ack_1 : boolean;
  signal ptr_deref_2829_store_0_req_0 : boolean;
  signal ptr_deref_2829_store_0_ack_0 : boolean;
  signal ptr_deref_2829_store_0_req_1 : boolean;
  signal ptr_deref_2829_store_0_ack_1 : boolean;
  signal type_cast_2834_inst_req_0 : boolean;
  signal type_cast_2834_inst_ack_0 : boolean;
  signal type_cast_2834_inst_req_1 : boolean;
  signal type_cast_2834_inst_ack_1 : boolean;
  signal if_stmt_2847_branch_req_0 : boolean;
  signal if_stmt_2847_branch_ack_1 : boolean;
  signal if_stmt_2847_branch_ack_0 : boolean;
  signal type_cast_2875_inst_req_0 : boolean;
  signal type_cast_2875_inst_ack_0 : boolean;
  signal type_cast_2875_inst_req_1 : boolean;
  signal type_cast_2875_inst_ack_1 : boolean;
  signal if_stmt_2894_branch_req_0 : boolean;
  signal if_stmt_2894_branch_ack_1 : boolean;
  signal if_stmt_2894_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2930_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2930_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2930_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2930_inst_ack_1 : boolean;
  signal phi_stmt_2697_req_0 : boolean;
  signal phi_stmt_2704_req_0 : boolean;
  signal phi_stmt_2711_req_0 : boolean;
  signal type_cast_2721_inst_req_0 : boolean;
  signal type_cast_2721_inst_ack_0 : boolean;
  signal type_cast_2721_inst_req_1 : boolean;
  signal type_cast_2721_inst_ack_1 : boolean;
  signal phi_stmt_2718_req_0 : boolean;
  signal type_cast_2703_inst_req_0 : boolean;
  signal type_cast_2703_inst_ack_0 : boolean;
  signal type_cast_2703_inst_req_1 : boolean;
  signal type_cast_2703_inst_ack_1 : boolean;
  signal phi_stmt_2697_req_1 : boolean;
  signal type_cast_2710_inst_req_0 : boolean;
  signal type_cast_2710_inst_ack_0 : boolean;
  signal type_cast_2710_inst_req_1 : boolean;
  signal type_cast_2710_inst_ack_1 : boolean;
  signal phi_stmt_2704_req_1 : boolean;
  signal type_cast_2717_inst_req_0 : boolean;
  signal type_cast_2717_inst_ack_0 : boolean;
  signal type_cast_2717_inst_req_1 : boolean;
  signal type_cast_2717_inst_ack_1 : boolean;
  signal phi_stmt_2711_req_1 : boolean;
  signal type_cast_2723_inst_req_0 : boolean;
  signal type_cast_2723_inst_ack_0 : boolean;
  signal type_cast_2723_inst_req_1 : boolean;
  signal type_cast_2723_inst_ack_1 : boolean;
  signal phi_stmt_2718_req_1 : boolean;
  signal phi_stmt_2697_ack_0 : boolean;
  signal phi_stmt_2704_ack_0 : boolean;
  signal phi_stmt_2711_ack_0 : boolean;
  signal phi_stmt_2718_ack_0 : boolean;
  signal phi_stmt_2901_req_1 : boolean;
  signal type_cast_2913_inst_req_0 : boolean;
  signal type_cast_2913_inst_ack_0 : boolean;
  signal type_cast_2913_inst_req_1 : boolean;
  signal type_cast_2913_inst_ack_1 : boolean;
  signal phi_stmt_2908_req_1 : boolean;
  signal type_cast_2919_inst_req_0 : boolean;
  signal type_cast_2919_inst_ack_0 : boolean;
  signal type_cast_2919_inst_req_1 : boolean;
  signal type_cast_2919_inst_ack_1 : boolean;
  signal phi_stmt_2914_req_1 : boolean;
  signal type_cast_2904_inst_req_0 : boolean;
  signal type_cast_2904_inst_ack_0 : boolean;
  signal type_cast_2904_inst_req_1 : boolean;
  signal type_cast_2904_inst_ack_1 : boolean;
  signal phi_stmt_2901_req_0 : boolean;
  signal type_cast_2911_inst_req_0 : boolean;
  signal type_cast_2911_inst_ack_0 : boolean;
  signal type_cast_2911_inst_req_1 : boolean;
  signal type_cast_2911_inst_ack_1 : boolean;
  signal phi_stmt_2908_req_0 : boolean;
  signal type_cast_2917_inst_req_0 : boolean;
  signal type_cast_2917_inst_ack_0 : boolean;
  signal type_cast_2917_inst_req_1 : boolean;
  signal type_cast_2917_inst_ack_1 : boolean;
  signal phi_stmt_2914_req_0 : boolean;
  signal phi_stmt_2901_ack_0 : boolean;
  signal phi_stmt_2908_ack_0 : boolean;
  signal phi_stmt_2914_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6778_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6778_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6778_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6778_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6778: Block -- control-path 
    signal convTransposeD_CP_6778_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6778_elements(0) <= convTransposeD_CP_6778_start;
    convTransposeD_CP_6778_symbol <= convTransposeD_CP_6778_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/$entry
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642__entry__
      -- CP-element group 0: 	 branch_block_stmt_2581/branch_block_stmt_2581__entry__
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2581/$entry
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_update_start_
      -- 
    cr_6999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(0), ack => type_cast_2627_inst_req_1); -- 
    rr_6826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(0), ack => RPIPE_Block3_start_2583_inst_req_0); -- 
    cr_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(0), ack => type_cast_2614_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2581/assign_stmt_2926__exit__
      -- CP-element group 1: 	 branch_block_stmt_2581/assign_stmt_2926__entry__
      -- CP-element group 1: 	 branch_block_stmt_2581/merge_stmt_2900__exit__
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2581/assign_stmt_2926/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/assign_stmt_2926/$exit
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/Update/cr
      -- 
    rr_7499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2703_inst_req_0); -- 
    cr_7504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2703_inst_req_1); -- 
    rr_7522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2710_inst_req_0); -- 
    cr_7527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2710_inst_req_1); -- 
    rr_7545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2717_inst_req_0); -- 
    cr_7550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2717_inst_req_1); -- 
    rr_7568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2723_inst_req_0); -- 
    cr_7573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(1), ack => type_cast_2723_inst_req_1); -- 
    convTransposeD_CP_6778_elements(1) <= convTransposeD_CP_6778_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_Sample/$exit
      -- 
    ra_6827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2583_inst_ack_0, ack => convTransposeD_CP_6778_elements(2)); -- 
    cr_6831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(2), ack => RPIPE_Block3_start_2583_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2583_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_Sample/rr
      -- 
    ca_6832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2583_inst_ack_1, ack => convTransposeD_CP_6778_elements(3)); -- 
    rr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(3), ack => RPIPE_Block3_start_2586_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_Sample/ra
      -- 
    ra_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2586_inst_ack_0, ack => convTransposeD_CP_6778_elements(4)); -- 
    cr_6845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(4), ack => RPIPE_Block3_start_2586_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2586_Update/ca
      -- 
    ca_6846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2586_inst_ack_1, ack => convTransposeD_CP_6778_elements(5)); -- 
    rr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(5), ack => RPIPE_Block3_start_2589_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_sample_completed_
      -- 
    ra_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2589_inst_ack_0, ack => convTransposeD_CP_6778_elements(6)); -- 
    cr_6859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(6), ack => RPIPE_Block3_start_2589_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2589_Update/ca
      -- 
    ca_6860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2589_inst_ack_1, ack => convTransposeD_CP_6778_elements(7)); -- 
    rr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(7), ack => RPIPE_Block3_start_2592_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_Update/cr
      -- 
    ra_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2592_inst_ack_0, ack => convTransposeD_CP_6778_elements(8)); -- 
    cr_6873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(8), ack => RPIPE_Block3_start_2592_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2592_Update/$exit
      -- 
    ca_6874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2592_inst_ack_1, ack => convTransposeD_CP_6778_elements(9)); -- 
    rr_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(9), ack => RPIPE_Block3_start_2595_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_Sample/ra
      -- 
    ra_6883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2595_inst_ack_0, ack => convTransposeD_CP_6778_elements(10)); -- 
    cr_6887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(10), ack => RPIPE_Block3_start_2595_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2595_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_Sample/rr
      -- 
    ca_6888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2595_inst_ack_1, ack => convTransposeD_CP_6778_elements(11)); -- 
    rr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(11), ack => RPIPE_Block3_start_2598_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_Sample/ra
      -- 
    ra_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2598_inst_ack_0, ack => convTransposeD_CP_6778_elements(12)); -- 
    cr_6901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(12), ack => RPIPE_Block3_start_2598_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2598_Update/$exit
      -- 
    ca_6902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2598_inst_ack_1, ack => convTransposeD_CP_6778_elements(13)); -- 
    rr_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(13), ack => RPIPE_Block3_start_2601_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_sample_completed_
      -- 
    ra_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2601_inst_ack_0, ack => convTransposeD_CP_6778_elements(14)); -- 
    cr_6915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(14), ack => RPIPE_Block3_start_2601_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2601_update_completed_
      -- 
    ca_6916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2601_inst_ack_1, ack => convTransposeD_CP_6778_elements(15)); -- 
    rr_6924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(15), ack => RPIPE_Block3_start_2604_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_Update/$entry
      -- 
    ra_6925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2604_inst_ack_0, ack => convTransposeD_CP_6778_elements(16)); -- 
    cr_6929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(16), ack => RPIPE_Block3_start_2604_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2604_Update/$exit
      -- 
    ca_6930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2604_inst_ack_1, ack => convTransposeD_CP_6778_elements(17)); -- 
    rr_6938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(17), ack => RPIPE_Block3_start_2607_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_update_start_
      -- 
    ra_6939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2607_inst_ack_0, ack => convTransposeD_CP_6778_elements(18)); -- 
    cr_6943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(18), ack => RPIPE_Block3_start_2607_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2607_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_sample_start_
      -- 
    ca_6944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2607_inst_ack_1, ack => convTransposeD_CP_6778_elements(19)); -- 
    rr_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(19), ack => RPIPE_Block3_start_2610_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_sample_completed_
      -- 
    ra_6953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2610_inst_ack_0, ack => convTransposeD_CP_6778_elements(20)); -- 
    cr_6957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(20), ack => RPIPE_Block3_start_2610_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2610_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_Sample/$entry
      -- 
    ca_6958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2610_inst_ack_1, ack => convTransposeD_CP_6778_elements(21)); -- 
    rr_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(21), ack => type_cast_2614_inst_req_0); -- 
    rr_6980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(21), ack => RPIPE_Block3_start_2623_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_sample_completed_
      -- 
    ra_6967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_0, ack => convTransposeD_CP_6778_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2614_Update/$exit
      -- 
    ca_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_1, ack => convTransposeD_CP_6778_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_update_start_
      -- 
    ra_6981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2623_inst_ack_0, ack => convTransposeD_CP_6778_elements(24)); -- 
    cr_6985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(24), ack => RPIPE_Block3_start_2623_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2623_update_completed_
      -- 
    ca_6986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2623_inst_ack_1, ack => convTransposeD_CP_6778_elements(25)); -- 
    rr_6994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(25), ack => type_cast_2627_inst_req_0); -- 
    rr_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(25), ack => RPIPE_Block3_start_2635_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_sample_completed_
      -- 
    ra_6995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2627_inst_ack_0, ack => convTransposeD_CP_6778_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/type_cast_2627_update_completed_
      -- 
    ca_7000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2627_inst_ack_1, ack => convTransposeD_CP_6778_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_Update/cr
      -- 
    ra_7009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2635_inst_ack_0, ack => convTransposeD_CP_6778_elements(28)); -- 
    cr_7013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(28), ack => RPIPE_Block3_start_2635_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2635_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_sample_start_
      -- 
    ca_7014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2635_inst_ack_1, ack => convTransposeD_CP_6778_elements(29)); -- 
    rr_7022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(29), ack => RPIPE_Block3_start_2638_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_sample_completed_
      -- 
    ra_7023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2638_inst_ack_0, ack => convTransposeD_CP_6778_elements(30)); -- 
    cr_7027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(30), ack => RPIPE_Block3_start_2638_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2638_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_sample_start_
      -- 
    ca_7028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2638_inst_ack_1, ack => convTransposeD_CP_6778_elements(31)); -- 
    rr_7036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(31), ack => RPIPE_Block3_start_2641_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_update_start_
      -- 
    ra_7037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2641_inst_ack_0, ack => convTransposeD_CP_6778_elements(32)); -- 
    cr_7041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(32), ack => RPIPE_Block3_start_2641_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/RPIPE_Block3_start_2641_Update/ca
      -- 
    ca_7042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2641_inst_ack_1, ack => convTransposeD_CP_6778_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/$entry
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642/$exit
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2584_to_assign_stmt_2642__exit__
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694__entry__
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_Sample/$entry
      -- 
    cr_7072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2689_inst_req_1); -- 
    cr_7086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2693_inst_req_1); -- 
    cr_7058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2685_inst_req_1); -- 
    rr_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2689_inst_req_0); -- 
    rr_7053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2685_inst_req_0); -- 
    rr_7081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(34), ack => type_cast_2693_inst_req_0); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(23) & convTransposeD_CP_6778_elements(27) & convTransposeD_CP_6778_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_Sample/ra
      -- 
    ra_7054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2685_inst_ack_0, ack => convTransposeD_CP_6778_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2685_Update/$exit
      -- 
    ca_7059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2685_inst_ack_1, ack => convTransposeD_CP_6778_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_sample_completed_
      -- 
    ra_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2689_inst_ack_0, ack => convTransposeD_CP_6778_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2689_update_completed_
      -- 
    ca_7073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2689_inst_ack_1, ack => convTransposeD_CP_6778_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_Sample/$exit
      -- 
    ra_7082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2693_inst_ack_0, ack => convTransposeD_CP_6778_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/type_cast_2693_Update/ca
      -- 
    ca_7087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2693_inst_ack_1, ack => convTransposeD_CP_6778_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694/$exit
      -- CP-element group 41: 	 branch_block_stmt_2581/assign_stmt_2649_to_assign_stmt_2694__exit__
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2697/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2704/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2711/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/Update/cr
      -- 
    rr_7473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(41), ack => type_cast_2721_inst_req_0); -- 
    cr_7478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(41), ack => type_cast_2721_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(36) & convTransposeD_CP_6778_elements(38) & convTransposeD_CP_6778_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_Sample/ra
      -- 
    ra_7099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2758_inst_ack_0, ack => convTransposeD_CP_6778_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_Update/$exit
      -- 
    ca_7104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2758_inst_ack_1, ack => convTransposeD_CP_6778_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_Sample/ra
      -- 
    ra_7113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2762_inst_ack_0, ack => convTransposeD_CP_6778_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_Update/$exit
      -- 
    ca_7118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2762_inst_ack_1, ack => convTransposeD_CP_6778_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_sample_completed_
      -- 
    ra_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_0, ack => convTransposeD_CP_6778_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_Update/ca
      -- 
    ca_7132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_1, ack => convTransposeD_CP_6778_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_sample_completed_
      -- 
    ra_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2796_inst_ack_0, ack => convTransposeD_CP_6778_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_index_scale_1/scale_rename_ack
      -- 
    ca_7146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2796_inst_ack_1, ack => convTransposeD_CP_6778_elements(49)); -- 
    req_7171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(49), ack => array_obj_ref_2802_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_Sample/$exit
      -- 
    ack_7172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2802_index_offset_ack_0, ack => convTransposeD_CP_6778_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_request/req
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_sample_start_
      -- 
    ack_7177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2802_index_offset_ack_1, ack => convTransposeD_CP_6778_elements(51)); -- 
    req_7186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(51), ack => addr_of_2803_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_request/ack
      -- CP-element group 52: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_sample_completed_
      -- 
    ack_7187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2803_final_reg_ack_0, ack => convTransposeD_CP_6778_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Sample/word_access_start/word_0/rr
      -- 
    ack_7192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2803_final_reg_ack_1, ack => convTransposeD_CP_6778_elements(53)); -- 
    rr_7225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(53), ack => ptr_deref_2807_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Sample/word_access_start/word_0/ra
      -- 
    ra_7226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2807_load_0_ack_0, ack => convTransposeD_CP_6778_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/ptr_deref_2807_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/ptr_deref_2807_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/ptr_deref_2807_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/ptr_deref_2807_Merge/merge_ack
      -- 
    ca_7237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2807_load_0_ack_1, ack => convTransposeD_CP_6778_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_Sample/req
      -- 
    req_7267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(56), ack => array_obj_ref_2825_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(43) & convTransposeD_CP_6778_elements(45) & convTransposeD_CP_6778_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_Sample/ack
      -- 
    ack_7268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2825_index_offset_ack_0, ack => convTransposeD_CP_6778_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_request/req
      -- 
    ack_7273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2825_index_offset_ack_1, ack => convTransposeD_CP_6778_elements(58)); -- 
    req_7282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(58), ack => addr_of_2826_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_request/ack
      -- 
    ack_7283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2826_final_reg_ack_0, ack => convTransposeD_CP_6778_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_word_addrgen/root_register_ack
      -- 
    ack_7288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2826_final_reg_ack_1, ack => convTransposeD_CP_6778_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/ptr_deref_2829_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/ptr_deref_2829_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/ptr_deref_2829_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/ptr_deref_2829_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/word_access_start/word_0/rr
      -- 
    rr_7326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(61), ack => ptr_deref_2829_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(55) & convTransposeD_CP_6778_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Sample/word_access_start/word_0/ra
      -- 
    ra_7327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2829_store_0_ack_0, ack => convTransposeD_CP_6778_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Update/word_access_complete/word_0/ca
      -- 
    ca_7338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2829_store_0_ack_1, ack => convTransposeD_CP_6778_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_Sample/ra
      -- 
    ra_7347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2834_inst_ack_0, ack => convTransposeD_CP_6778_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_Update/ca
      -- 
    ca_7352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2834_inst_ack_1, ack => convTransposeD_CP_6778_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/$exit
      -- CP-element group 66: 	 branch_block_stmt_2581/if_stmt_2847__entry__
      -- CP-element group 66: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846__exit__
      -- CP-element group 66: 	 branch_block_stmt_2581/if_stmt_2847_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2581/if_stmt_2847_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2581/if_stmt_2847_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2581/if_stmt_2847_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2581/R_cmp_2848_place
      -- CP-element group 66: 	 branch_block_stmt_2581/if_stmt_2847_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2581/if_stmt_2847_else_link/$entry
      -- 
    branch_req_7360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(66), ack => if_stmt_2847_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(50) & convTransposeD_CP_6778_elements(57) & convTransposeD_CP_6778_elements(63) & convTransposeD_CP_6778_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2581/assign_stmt_2859__entry__
      -- CP-element group 67: 	 branch_block_stmt_2581/assign_stmt_2859__exit__
      -- CP-element group 67: 	 branch_block_stmt_2581/merge_stmt_2853__exit__
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2581/if_stmt_2847_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2581/if_stmt_2847_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2581/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2581/assign_stmt_2859/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/assign_stmt_2859/$exit
      -- CP-element group 67: 	 branch_block_stmt_2581/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2581/merge_stmt_2853_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2581/merge_stmt_2853_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/merge_stmt_2853_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2581/merge_stmt_2853_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2847_branch_ack_1, ack => convTransposeD_CP_6778_elements(67)); -- 
    rr_7683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2904_inst_req_0); -- 
    cr_7688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2904_inst_req_1); -- 
    rr_7706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2911_inst_req_0); -- 
    cr_7711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2911_inst_req_1); -- 
    rr_7729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2917_inst_req_0); -- 
    cr_7734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(67), ack => type_cast_2917_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893__entry__
      -- CP-element group 68: 	 branch_block_stmt_2581/merge_stmt_2861__exit__
      -- CP-element group 68: 	 branch_block_stmt_2581/if_stmt_2847_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2581/if_stmt_2847_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2581/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/$entry
      -- CP-element group 68: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2581/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2581/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2581/merge_stmt_2861_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2581/merge_stmt_2861_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2581/merge_stmt_2861_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2581/merge_stmt_2861_PhiAck/dummy
      -- 
    else_choice_transition_7369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2847_branch_ack_0, ack => convTransposeD_CP_6778_elements(68)); -- 
    rr_7385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(68), ack => type_cast_2875_inst_req_0); -- 
    cr_7390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(68), ack => type_cast_2875_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_Sample/ra
      -- 
    ra_7386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2875_inst_ack_0, ack => convTransposeD_CP_6778_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893__exit__
      -- CP-element group 70: 	 branch_block_stmt_2581/if_stmt_2894__entry__
      -- CP-element group 70: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/$exit
      -- CP-element group 70: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2581/assign_stmt_2867_to_assign_stmt_2893/type_cast_2875_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2581/if_stmt_2894_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2581/if_stmt_2894_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2581/if_stmt_2894_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2581/if_stmt_2894_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2581/R_cmp121_2895_place
      -- CP-element group 70: 	 branch_block_stmt_2581/if_stmt_2894_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2581/if_stmt_2894_else_link/$entry
      -- 
    ca_7391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2875_inst_ack_1, ack => convTransposeD_CP_6778_elements(70)); -- 
    branch_req_7399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(70), ack => if_stmt_2894_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2581/merge_stmt_2928__exit__
      -- CP-element group 71: 	 branch_block_stmt_2581/assign_stmt_2933__entry__
      -- CP-element group 71: 	 branch_block_stmt_2581/if_stmt_2894_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2581/if_stmt_2894_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2581/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2581/assign_stmt_2933/$entry
      -- CP-element group 71: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2581/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2581/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2581/merge_stmt_2928_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2581/merge_stmt_2928_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2581/merge_stmt_2928_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2581/merge_stmt_2928_PhiAck/dummy
      -- 
    if_choice_transition_7404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2894_branch_ack_1, ack => convTransposeD_CP_6778_elements(71)); -- 
    req_7424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(71), ack => WPIPE_Block3_done_2930_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2581/if_stmt_2894_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2581/if_stmt_2894_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2901/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2894_branch_ack_0, ack => convTransposeD_CP_6778_elements(72)); -- 
    rr_7634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(72), ack => type_cast_2913_inst_req_0); -- 
    cr_7639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(72), ack => type_cast_2913_inst_req_1); -- 
    rr_7657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(72), ack => type_cast_2919_inst_req_0); -- 
    cr_7662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(72), ack => type_cast_2919_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_Update/req
      -- 
    ack_7425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2930_inst_ack_0, ack => convTransposeD_CP_6778_elements(73)); -- 
    req_7429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(73), ack => WPIPE_Block3_done_2930_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 branch_block_stmt_2581/return__
      -- CP-element group 74: 	 branch_block_stmt_2581/merge_stmt_2935__exit__
      -- CP-element group 74: 	 branch_block_stmt_2581/branch_block_stmt_2581__exit__
      -- CP-element group 74: 	 branch_block_stmt_2581/$exit
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2581/assign_stmt_2933__exit__
      -- CP-element group 74: 	 branch_block_stmt_2581/assign_stmt_2933/$exit
      -- CP-element group 74: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2581/assign_stmt_2933/WPIPE_Block3_done_2930_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2581/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2581/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2581/merge_stmt_2935_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2581/merge_stmt_2935_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2581/merge_stmt_2935_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2581/merge_stmt_2935_PhiAck/dummy
      -- 
    ack_7430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2930_inst_ack_1, ack => convTransposeD_CP_6778_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2697/$exit
      -- CP-element group 75: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2701_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_req
      -- 
    phi_stmt_2697_req_7441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2697_req_7441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(75), ack => phi_stmt_2697_req_0); -- 
    -- Element group convTransposeD_CP_6778_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6778_elements(41), ack => convTransposeD_CP_6778_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2704/$exit
      -- CP-element group 76: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2708_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_req
      -- 
    phi_stmt_2704_req_7449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2704_req_7449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(76), ack => phi_stmt_2704_req_0); -- 
    -- Element group convTransposeD_CP_6778_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6778_elements(41), ack => convTransposeD_CP_6778_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2711/$exit
      -- CP-element group 77: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2715_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_req
      -- 
    phi_stmt_2711_req_7457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2711_req_7457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(77), ack => phi_stmt_2711_req_0); -- 
    -- Element group convTransposeD_CP_6778_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6778_elements(41), ack => convTransposeD_CP_6778_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/Sample/ra
      -- 
    ra_7474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_0, ack => convTransposeD_CP_6778_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/Update/ca
      -- 
    ca_7479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_1, ack => convTransposeD_CP_6778_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/$exit
      -- CP-element group 80: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/$exit
      -- CP-element group 80: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2721/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_req
      -- 
    phi_stmt_2718_req_7480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2718_req_7480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(80), ack => phi_stmt_2718_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(78) & convTransposeD_CP_6778_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2581/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(75) & convTransposeD_CP_6778_elements(76) & convTransposeD_CP_6778_elements(77) & convTransposeD_CP_6778_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/Sample/ra
      -- 
    ra_7500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2703_inst_ack_0, ack => convTransposeD_CP_6778_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/Update/ca
      -- 
    ca_7505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2703_inst_ack_1, ack => convTransposeD_CP_6778_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/$exit
      -- CP-element group 84: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/$exit
      -- CP-element group 84: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_sources/type_cast_2703/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2697/phi_stmt_2697_req
      -- 
    phi_stmt_2697_req_7506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2697_req_7506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(84), ack => phi_stmt_2697_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(82) & convTransposeD_CP_6778_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/Sample/ra
      -- 
    ra_7523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_0, ack => convTransposeD_CP_6778_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/Update/ca
      -- 
    ca_7528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_1, ack => convTransposeD_CP_6778_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/$exit
      -- CP-element group 87: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/$exit
      -- CP-element group 87: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_sources/type_cast_2710/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2704/phi_stmt_2704_req
      -- 
    phi_stmt_2704_req_7529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2704_req_7529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(87), ack => phi_stmt_2704_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(85) & convTransposeD_CP_6778_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/Sample/ra
      -- 
    ra_7546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2717_inst_ack_0, ack => convTransposeD_CP_6778_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/Update/ca
      -- 
    ca_7551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2717_inst_ack_1, ack => convTransposeD_CP_6778_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/$exit
      -- CP-element group 90: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/$exit
      -- CP-element group 90: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_sources/type_cast_2717/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2711/phi_stmt_2711_req
      -- 
    phi_stmt_2711_req_7552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2711_req_7552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(90), ack => phi_stmt_2711_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(88) & convTransposeD_CP_6778_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/Sample/ra
      -- 
    ra_7569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2723_inst_ack_0, ack => convTransposeD_CP_6778_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/Update/ca
      -- 
    ca_7574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2723_inst_ack_1, ack => convTransposeD_CP_6778_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/$exit
      -- CP-element group 93: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/$exit
      -- CP-element group 93: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_sources/type_cast_2723/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2718/phi_stmt_2718_req
      -- 
    phi_stmt_2718_req_7575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2718_req_7575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(93), ack => phi_stmt_2718_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(91) & convTransposeD_CP_6778_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2581/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(84) & convTransposeD_CP_6778_elements(87) & convTransposeD_CP_6778_elements(90) & convTransposeD_CP_6778_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2581/merge_stmt_2696_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2581/merge_stmt_2696_PhiAck/$entry
      -- 
    convTransposeD_CP_6778_elements(95) <= OrReduce(convTransposeD_CP_6778_elements(81) & convTransposeD_CP_6778_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2581/merge_stmt_2696_PhiAck/phi_stmt_2697_ack
      -- 
    phi_stmt_2697_ack_7580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2697_ack_0, ack => convTransposeD_CP_6778_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2581/merge_stmt_2696_PhiAck/phi_stmt_2704_ack
      -- 
    phi_stmt_2704_ack_7581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2704_ack_0, ack => convTransposeD_CP_6778_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2581/merge_stmt_2696_PhiAck/phi_stmt_2711_ack
      -- 
    phi_stmt_2711_ack_7582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2711_ack_0, ack => convTransposeD_CP_6778_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2581/merge_stmt_2696_PhiAck/phi_stmt_2718_ack
      -- 
    phi_stmt_2718_ack_7583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2718_ack_0, ack => convTransposeD_CP_6778_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/merge_stmt_2696__exit__
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846__entry__
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2758_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2803_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2796_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2802_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2762_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2766_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2807_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/array_obj_ref_2825_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/addr_of_2826_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/ptr_deref_2829_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2581/assign_stmt_2730_to_assign_stmt_2846/type_cast_2834_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2581/merge_stmt_2696_PhiAck/$exit
      -- 
    rr_7098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2758_inst_req_0); -- 
    cr_7103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2758_inst_req_1); -- 
    cr_7117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2762_inst_req_1); -- 
    rr_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2766_inst_req_0); -- 
    rr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2796_inst_req_0); -- 
    cr_7145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2796_inst_req_1); -- 
    req_7191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => addr_of_2803_final_reg_req_1); -- 
    req_7176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => array_obj_ref_2802_index_offset_req_1); -- 
    cr_7131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2766_inst_req_1); -- 
    rr_7112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2762_inst_req_0); -- 
    cr_7236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => ptr_deref_2807_load_0_req_1); -- 
    req_7272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => array_obj_ref_2825_index_offset_req_1); -- 
    req_7287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => addr_of_2826_final_reg_req_1); -- 
    cr_7337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => ptr_deref_2829_store_0_req_1); -- 
    rr_7346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2834_inst_req_0); -- 
    cr_7351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(100), ack => type_cast_2834_inst_req_1); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(96) & convTransposeD_CP_6778_elements(97) & convTransposeD_CP_6778_elements(98) & convTransposeD_CP_6778_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2901/$exit
      -- CP-element group 101: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2907_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_req
      -- 
    phi_stmt_2901_req_7618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2901_req_7618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(101), ack => phi_stmt_2901_req_1); -- 
    -- Element group convTransposeD_CP_6778_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6778_elements(72), ack => convTransposeD_CP_6778_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Sample/ra
      -- 
    ra_7635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2913_inst_ack_0, ack => convTransposeD_CP_6778_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/Update/ca
      -- 
    ca_7640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2913_inst_ack_1, ack => convTransposeD_CP_6778_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/$exit
      -- CP-element group 104: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/$exit
      -- CP-element group 104: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2913/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_req
      -- 
    phi_stmt_2908_req_7641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2908_req_7641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(104), ack => phi_stmt_2908_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(102) & convTransposeD_CP_6778_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Sample/ra
      -- 
    ra_7658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2919_inst_ack_0, ack => convTransposeD_CP_6778_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/Update/ca
      -- 
    ca_7663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2919_inst_ack_1, ack => convTransposeD_CP_6778_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/$exit
      -- CP-element group 107: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/$exit
      -- CP-element group 107: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2919/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_req
      -- 
    phi_stmt_2914_req_7664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2914_req_7664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(107), ack => phi_stmt_2914_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(105) & convTransposeD_CP_6778_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2581/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(101) & convTransposeD_CP_6778_elements(104) & convTransposeD_CP_6778_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/Sample/ra
      -- 
    ra_7684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2904_inst_ack_0, ack => convTransposeD_CP_6778_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/Update/ca
      -- 
    ca_7689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2904_inst_ack_1, ack => convTransposeD_CP_6778_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/$exit
      -- CP-element group 111: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/$exit
      -- CP-element group 111: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_sources/type_cast_2904/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2901/phi_stmt_2901_req
      -- 
    phi_stmt_2901_req_7690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2901_req_7690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(111), ack => phi_stmt_2901_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(109) & convTransposeD_CP_6778_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Sample/ra
      -- 
    ra_7707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2911_inst_ack_0, ack => convTransposeD_CP_6778_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/Update/ca
      -- 
    ca_7712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2911_inst_ack_1, ack => convTransposeD_CP_6778_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/$exit
      -- CP-element group 114: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/$exit
      -- CP-element group 114: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_sources/type_cast_2911/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2908/phi_stmt_2908_req
      -- 
    phi_stmt_2908_req_7713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2908_req_7713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(114), ack => phi_stmt_2908_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(112) & convTransposeD_CP_6778_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Sample/ra
      -- 
    ra_7730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2917_inst_ack_0, ack => convTransposeD_CP_6778_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/Update/ca
      -- 
    ca_7735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2917_inst_ack_1, ack => convTransposeD_CP_6778_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/$exit
      -- CP-element group 117: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/$exit
      -- CP-element group 117: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_sources/type_cast_2917/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2914/phi_stmt_2914_req
      -- 
    phi_stmt_2914_req_7736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2914_req_7736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6778_elements(117), ack => phi_stmt_2914_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(115) & convTransposeD_CP_6778_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2581/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(111) & convTransposeD_CP_6778_elements(114) & convTransposeD_CP_6778_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2581/merge_stmt_2900_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2581/merge_stmt_2900_PhiAck/$entry
      -- 
    convTransposeD_CP_6778_elements(119) <= OrReduce(convTransposeD_CP_6778_elements(108) & convTransposeD_CP_6778_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2581/merge_stmt_2900_PhiAck/phi_stmt_2901_ack
      -- 
    phi_stmt_2901_ack_7741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2901_ack_0, ack => convTransposeD_CP_6778_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2581/merge_stmt_2900_PhiAck/phi_stmt_2908_ack
      -- 
    phi_stmt_2908_ack_7742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2908_ack_0, ack => convTransposeD_CP_6778_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2581/merge_stmt_2900_PhiAck/phi_stmt_2914_ack
      -- 
    phi_stmt_2914_ack_7743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2914_ack_0, ack => convTransposeD_CP_6778_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2581/merge_stmt_2900_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6778_elements(120) & convTransposeD_CP_6778_elements(121) & convTransposeD_CP_6778_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6778_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2824_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2824_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2801_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2801_scaled : std_logic_vector(13 downto 0);
    signal add103_2859 : std_logic_vector(15 downto 0);
    signal add32_2660 : std_logic_vector(15 downto 0);
    signal add50_2666 : std_logic_vector(15 downto 0);
    signal add63_2677 : std_logic_vector(15 downto 0);
    signal add82_2777 : std_logic_vector(63 downto 0);
    signal add84_2787 : std_logic_vector(63 downto 0);
    signal add96_2841 : std_logic_vector(31 downto 0);
    signal add_2633 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2735 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2802_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2802_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2802_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2802_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2802_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2802_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2825_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2825_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2825_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2825_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2825_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2825_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2804 : std_logic_vector(31 downto 0);
    signal arrayidx92_2827 : std_logic_vector(31 downto 0);
    signal call11_2602 : std_logic_vector(15 downto 0);
    signal call13_2605 : std_logic_vector(15 downto 0);
    signal call14_2608 : std_logic_vector(15 downto 0);
    signal call15_2611 : std_logic_vector(15 downto 0);
    signal call16_2624 : std_logic_vector(15 downto 0);
    signal call18_2636 : std_logic_vector(15 downto 0);
    signal call1_2587 : std_logic_vector(15 downto 0);
    signal call20_2639 : std_logic_vector(15 downto 0);
    signal call22_2642 : std_logic_vector(15 downto 0);
    signal call3_2590 : std_logic_vector(15 downto 0);
    signal call5_2593 : std_logic_vector(15 downto 0);
    signal call7_2596 : std_logic_vector(15 downto 0);
    signal call9_2599 : std_logic_vector(15 downto 0);
    signal call_2584 : std_logic_vector(15 downto 0);
    signal cmp111_2872 : std_logic_vector(0 downto 0);
    signal cmp121_2893 : std_logic_vector(0 downto 0);
    signal cmp_2846 : std_logic_vector(0 downto 0);
    signal conv17_2628 : std_logic_vector(31 downto 0);
    signal conv70_2759 : std_logic_vector(63 downto 0);
    signal conv73_2686 : std_logic_vector(63 downto 0);
    signal conv75_2763 : std_logic_vector(63 downto 0);
    signal conv78_2690 : std_logic_vector(63 downto 0);
    signal conv80_2767 : std_logic_vector(63 downto 0);
    signal conv95_2835 : std_logic_vector(31 downto 0);
    signal conv99_2694 : std_logic_vector(31 downto 0);
    signal conv_2615 : std_logic_vector(31 downto 0);
    signal idxprom91_2820 : std_logic_vector(63 downto 0);
    signal idxprom_2797 : std_logic_vector(63 downto 0);
    signal inc115_2876 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2881 : std_logic_vector(15 downto 0);
    signal inc_2867 : std_logic_vector(15 downto 0);
    signal indvar_2697 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2926 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2914 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2718 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2908 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2711 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2888 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2901 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2704 : std_logic_vector(15 downto 0);
    signal mul59_2750 : std_logic_vector(15 downto 0);
    signal mul81_2772 : std_logic_vector(63 downto 0);
    signal mul83_2782 : std_logic_vector(63 downto 0);
    signal mul_2740 : std_logic_vector(15 downto 0);
    signal ptr_deref_2807_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2807_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2807_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2807_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2807_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2829_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2829_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2829_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2829_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2829_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2829_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2621 : std_logic_vector(31 downto 0);
    signal shr135_2649 : std_logic_vector(15 downto 0);
    signal shr31136_2655 : std_logic_vector(15 downto 0);
    signal shr86_2793 : std_logic_vector(31 downto 0);
    signal shr90_2814 : std_logic_vector(63 downto 0);
    signal sub53_2745 : std_logic_vector(15 downto 0);
    signal sub66_2682 : std_logic_vector(15 downto 0);
    signal sub67_2755 : std_logic_vector(15 downto 0);
    signal sub_2671 : std_logic_vector(15 downto 0);
    signal tmp1_2730 : std_logic_vector(31 downto 0);
    signal tmp88_2808 : std_logic_vector(63 downto 0);
    signal type_cast_2619_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2647_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2653_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2664_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2675_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2701_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2703_wire : std_logic_vector(31 downto 0);
    signal type_cast_2708_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2710_wire : std_logic_vector(15 downto 0);
    signal type_cast_2715_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2717_wire : std_logic_vector(15 downto 0);
    signal type_cast_2721_wire : std_logic_vector(15 downto 0);
    signal type_cast_2723_wire : std_logic_vector(15 downto 0);
    signal type_cast_2728_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2791_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2812_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2818_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2839_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2857_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2865_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2885_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2904_wire : std_logic_vector(15 downto 0);
    signal type_cast_2907_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2911_wire : std_logic_vector(15 downto 0);
    signal type_cast_2913_wire : std_logic_vector(15 downto 0);
    signal type_cast_2917_wire : std_logic_vector(15 downto 0);
    signal type_cast_2919_wire : std_logic_vector(15 downto 0);
    signal type_cast_2924_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2932_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2802_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2802_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2802_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2802_resized_base_address <= "00000000000000";
    array_obj_ref_2825_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2825_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2825_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2825_resized_base_address <= "00000000000000";
    ptr_deref_2807_word_offset_0 <= "00000000000000";
    ptr_deref_2829_word_offset_0 <= "00000000000000";
    type_cast_2619_wire_constant <= "00000000000000000000000000010000";
    type_cast_2647_wire_constant <= "0000000000000010";
    type_cast_2653_wire_constant <= "0000000000000001";
    type_cast_2664_wire_constant <= "1111111111111111";
    type_cast_2675_wire_constant <= "1111111111111111";
    type_cast_2701_wire_constant <= "00000000000000000000000000000000";
    type_cast_2708_wire_constant <= "0000000000000000";
    type_cast_2715_wire_constant <= "0000000000000000";
    type_cast_2728_wire_constant <= "00000000000000000000000000000100";
    type_cast_2791_wire_constant <= "00000000000000000000000000000010";
    type_cast_2812_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2818_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2839_wire_constant <= "00000000000000000000000000000100";
    type_cast_2857_wire_constant <= "0000000000000100";
    type_cast_2865_wire_constant <= "0000000000000001";
    type_cast_2885_wire_constant <= "0000000000000000";
    type_cast_2907_wire_constant <= "0000000000000000";
    type_cast_2924_wire_constant <= "00000000000000000000000000000001";
    type_cast_2932_wire_constant <= "0000000000000001";
    phi_stmt_2697: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2701_wire_constant & type_cast_2703_wire;
      req <= phi_stmt_2697_req_0 & phi_stmt_2697_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2697",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2697_ack_0,
          idata => idata,
          odata => indvar_2697,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2697
    phi_stmt_2704: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2708_wire_constant & type_cast_2710_wire;
      req <= phi_stmt_2704_req_0 & phi_stmt_2704_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2704",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2704_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2704,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2704
    phi_stmt_2711: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2715_wire_constant & type_cast_2717_wire;
      req <= phi_stmt_2711_req_0 & phi_stmt_2711_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2711",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2711_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2711,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2711
    phi_stmt_2718: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2721_wire & type_cast_2723_wire;
      req <= phi_stmt_2718_req_0 & phi_stmt_2718_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2718",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2718_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2718,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2718
    phi_stmt_2901: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2904_wire & type_cast_2907_wire_constant;
      req <= phi_stmt_2901_req_0 & phi_stmt_2901_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2901",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2901_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2901,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2901
    phi_stmt_2908: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2911_wire & type_cast_2913_wire;
      req <= phi_stmt_2908_req_0 & phi_stmt_2908_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2908",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2908_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2908,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2908
    phi_stmt_2914: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2917_wire & type_cast_2919_wire;
      req <= phi_stmt_2914_req_0 & phi_stmt_2914_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2914",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2914_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2914,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2914
    -- flow-through select operator MUX_2887_inst
    input_dim1x_x2_2888 <= type_cast_2885_wire_constant when (cmp111_2872(0) /=  '0') else inc_2867;
    addr_of_2803_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2803_final_reg_req_0;
      addr_of_2803_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2803_final_reg_req_1;
      addr_of_2803_final_reg_ack_1<= rack(0);
      addr_of_2803_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2803_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2802_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2804,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2826_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2826_final_reg_req_0;
      addr_of_2826_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2826_final_reg_req_1;
      addr_of_2826_final_reg_ack_1<= rack(0);
      addr_of_2826_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2826_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2825_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2827,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2614_inst_req_0;
      type_cast_2614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2614_inst_req_1;
      type_cast_2614_inst_ack_1<= rack(0);
      type_cast_2614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2627_inst_req_0;
      type_cast_2627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2627_inst_req_1;
      type_cast_2627_inst_ack_1<= rack(0);
      type_cast_2627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2624,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2628,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2685_inst_req_0;
      type_cast_2685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2685_inst_req_1;
      type_cast_2685_inst_ack_1<= rack(0);
      type_cast_2685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2642,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2689_inst_req_0;
      type_cast_2689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2689_inst_req_1;
      type_cast_2689_inst_ack_1<= rack(0);
      type_cast_2689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2639,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2693_inst_req_0;
      type_cast_2693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2693_inst_req_1;
      type_cast_2693_inst_ack_1<= rack(0);
      type_cast_2693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2694,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2703_inst_req_0;
      type_cast_2703_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2703_inst_req_1;
      type_cast_2703_inst_ack_1<= rack(0);
      type_cast_2703_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2703_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2926,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2703_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2710_inst_req_0;
      type_cast_2710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2710_inst_req_1;
      type_cast_2710_inst_ack_1<= rack(0);
      type_cast_2710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2710_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2717_inst_req_0;
      type_cast_2717_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2717_inst_req_1;
      type_cast_2717_inst_ack_1<= rack(0);
      type_cast_2717_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2717_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2717_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2721_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2721_inst_req_0;
      type_cast_2721_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2721_inst_req_1;
      type_cast_2721_inst_ack_1<= rack(0);
      type_cast_2721_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2721_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2721_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2723_inst_req_0;
      type_cast_2723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2723_inst_req_1;
      type_cast_2723_inst_ack_1<= rack(0);
      type_cast_2723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2914,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2723_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2758_inst_req_0;
      type_cast_2758_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2758_inst_req_1;
      type_cast_2758_inst_ack_1<= rack(0);
      type_cast_2758_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2758_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2704,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2759,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2762_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2762_inst_req_0;
      type_cast_2762_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2762_inst_req_1;
      type_cast_2762_inst_ack_1<= rack(0);
      type_cast_2762_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2762_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2763,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2766_inst_req_0;
      type_cast_2766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2766_inst_req_1;
      type_cast_2766_inst_ack_1<= rack(0);
      type_cast_2766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2745,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2767,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2796_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2796_inst_req_0;
      type_cast_2796_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2796_inst_req_1;
      type_cast_2796_inst_ack_1<= rack(0);
      type_cast_2796_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2796_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2793,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2834_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2834_inst_req_0;
      type_cast_2834_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2834_inst_req_1;
      type_cast_2834_inst_ack_1<= rack(0);
      type_cast_2834_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2834_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2704,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2835,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2875_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2875_inst_req_0;
      type_cast_2875_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2875_inst_req_1;
      type_cast_2875_inst_ack_1<= rack(0);
      type_cast_2875_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2875_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2876,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2904_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2904_inst_req_0;
      type_cast_2904_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2904_inst_req_1;
      type_cast_2904_inst_ack_1<= rack(0);
      type_cast_2904_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2904_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2859,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2904_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2911_inst_req_0;
      type_cast_2911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2911_inst_req_1;
      type_cast_2911_inst_ack_1<= rack(0);
      type_cast_2911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2911_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2711,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2911_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2913_inst_req_0;
      type_cast_2913_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2913_inst_req_1;
      type_cast_2913_inst_ack_1<= rack(0);
      type_cast_2913_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2913_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2888,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2913_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2917_inst_req_0;
      type_cast_2917_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2917_inst_req_1;
      type_cast_2917_inst_ack_1<= rack(0);
      type_cast_2917_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2718,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2917_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2919_inst_req_0;
      type_cast_2919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2919_inst_req_1;
      type_cast_2919_inst_ack_1<= rack(0);
      type_cast_2919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2881,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2919_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2802_index_1_rename
    process(R_idxprom_2801_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2801_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2801_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2802_index_1_resize
    process(idxprom_2797) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2797;
      ov := iv(13 downto 0);
      R_idxprom_2801_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2802_root_address_inst
    process(array_obj_ref_2802_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2802_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2802_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2825_index_1_rename
    process(R_idxprom91_2824_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2824_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2824_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2825_index_1_resize
    process(idxprom91_2820) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2820;
      ov := iv(13 downto 0);
      R_idxprom91_2824_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2825_root_address_inst
    process(array_obj_ref_2825_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2825_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2825_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2807_addr_0
    process(ptr_deref_2807_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2807_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2807_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2807_base_resize
    process(arrayidx87_2804) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2804;
      ov := iv(13 downto 0);
      ptr_deref_2807_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2807_gather_scatter
    process(ptr_deref_2807_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2807_data_0;
      ov(63 downto 0) := iv;
      tmp88_2808 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2807_root_address_inst
    process(ptr_deref_2807_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2807_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2807_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2829_addr_0
    process(ptr_deref_2829_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2829_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2829_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2829_base_resize
    process(arrayidx92_2827) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2827;
      ov := iv(13 downto 0);
      ptr_deref_2829_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2829_gather_scatter
    process(tmp88_2808) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2808;
      ov(63 downto 0) := iv;
      ptr_deref_2829_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2829_root_address_inst
    process(ptr_deref_2829_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2829_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2829_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2847_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2846;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2847_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2847_branch_req_0,
          ack0 => if_stmt_2847_branch_ack_0,
          ack1 => if_stmt_2847_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2894_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2893;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2894_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2894_branch_req_0,
          ack0 => if_stmt_2894_branch_ack_0,
          ack1 => if_stmt_2894_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2659_inst
    process(shr135_2649, shr31136_2655) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2649, shr31136_2655, tmp_var);
      add32_2660 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2665_inst
    process(call7_2596) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2596, type_cast_2664_wire_constant, tmp_var);
      add50_2666 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2676_inst
    process(call9_2599) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2599, type_cast_2675_wire_constant, tmp_var);
      add63_2677 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2744_inst
    process(sub_2671, mul_2740) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2671, mul_2740, tmp_var);
      sub53_2745 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2754_inst
    process(sub66_2682, mul59_2750) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2682, mul59_2750, tmp_var);
      sub67_2755 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2858_inst
    process(input_dim2x_x1_2704) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2704, type_cast_2857_wire_constant, tmp_var);
      add103_2859 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2866_inst
    process(input_dim1x_x1_2711) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2711, type_cast_2865_wire_constant, tmp_var);
      inc_2867 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2880_inst
    process(inc115_2876, input_dim0x_x2_2718) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2876, input_dim0x_x2_2718, tmp_var);
      inc115x_xinput_dim0x_x2_2881 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2734_inst
    process(add_2633, tmp1_2730) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2633, tmp1_2730, tmp_var);
      add_src_0x_x0_2735 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2840_inst
    process(conv95_2835) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2835, type_cast_2839_wire_constant, tmp_var);
      add96_2841 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2925_inst
    process(indvar_2697) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2697, type_cast_2924_wire_constant, tmp_var);
      indvarx_xnext_2926 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2776_inst
    process(mul81_2772, conv75_2763) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2772, conv75_2763, tmp_var);
      add82_2777 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2786_inst
    process(mul83_2782, conv70_2759) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2782, conv70_2759, tmp_var);
      add84_2787 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2819_inst
    process(shr90_2814) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2814, type_cast_2818_wire_constant, tmp_var);
      idxprom91_2820 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2871_inst
    process(inc_2867, call1_2587) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2867, call1_2587, tmp_var);
      cmp111_2872 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2892_inst
    process(inc115x_xinput_dim0x_x2_2881, call_2584) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2881, call_2584, tmp_var);
      cmp121_2893 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2648_inst
    process(call_2584) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2584, type_cast_2647_wire_constant, tmp_var);
      shr135_2649 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2654_inst
    process(call_2584) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2584, type_cast_2653_wire_constant, tmp_var);
      shr31136_2655 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2792_inst
    process(add_src_0x_x0_2735) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2735, type_cast_2791_wire_constant, tmp_var);
      shr86_2793 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2813_inst
    process(add84_2787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2787, type_cast_2812_wire_constant, tmp_var);
      shr90_2814 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2739_inst
    process(input_dim0x_x2_2718, call13_2605) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2718, call13_2605, tmp_var);
      mul_2740 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2749_inst
    process(input_dim1x_x1_2711, call13_2605) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2711, call13_2605, tmp_var);
      mul59_2750 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2729_inst
    process(indvar_2697) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2697, type_cast_2728_wire_constant, tmp_var);
      tmp1_2730 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2771_inst
    process(conv80_2767, conv78_2690) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2767, conv78_2690, tmp_var);
      mul81_2772 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2781_inst
    process(add82_2777, conv73_2686) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2777, conv73_2686, tmp_var);
      mul83_2782 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2632_inst
    process(shl_2621, conv17_2628) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2621, conv17_2628, tmp_var);
      add_2633 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2620_inst
    process(conv_2615) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2615, type_cast_2619_wire_constant, tmp_var);
      shl_2621 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2670_inst
    process(add50_2666, call14_2608) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2666, call14_2608, tmp_var);
      sub_2671 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2681_inst
    process(add63_2677, call14_2608) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2677, call14_2608, tmp_var);
      sub66_2682 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2845_inst
    process(add96_2841, conv99_2694) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2841, conv99_2694, tmp_var);
      cmp_2846 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2802_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2801_scaled;
      array_obj_ref_2802_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2802_index_offset_req_0;
      array_obj_ref_2802_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2802_index_offset_req_1;
      array_obj_ref_2802_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2825_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2824_scaled;
      array_obj_ref_2825_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2825_index_offset_req_0;
      array_obj_ref_2825_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2825_index_offset_req_1;
      array_obj_ref_2825_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2807_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2807_load_0_req_0;
      ptr_deref_2807_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2807_load_0_req_1;
      ptr_deref_2807_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2807_word_address_0;
      ptr_deref_2807_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2829_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2829_store_0_req_0;
      ptr_deref_2829_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2829_store_0_req_1;
      ptr_deref_2829_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2829_word_address_0;
      data_in <= ptr_deref_2829_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2583_inst RPIPE_Block3_start_2586_inst RPIPE_Block3_start_2589_inst RPIPE_Block3_start_2592_inst RPIPE_Block3_start_2595_inst RPIPE_Block3_start_2598_inst RPIPE_Block3_start_2601_inst RPIPE_Block3_start_2604_inst RPIPE_Block3_start_2607_inst RPIPE_Block3_start_2610_inst RPIPE_Block3_start_2623_inst RPIPE_Block3_start_2635_inst RPIPE_Block3_start_2638_inst RPIPE_Block3_start_2641_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2583_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2586_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2589_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2592_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2595_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2598_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2601_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2604_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2607_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2610_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2623_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2635_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2638_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2641_inst_req_0;
      RPIPE_Block3_start_2583_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2586_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2589_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2592_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2595_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2598_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2601_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2604_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2607_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2610_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2623_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2635_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2638_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2641_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2583_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2586_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2589_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2592_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2595_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2598_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2601_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2604_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2607_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2610_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2623_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2635_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2638_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2641_inst_req_1;
      RPIPE_Block3_start_2583_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2586_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2589_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2592_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2595_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2598_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2601_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2604_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2607_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2610_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2623_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2635_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2638_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2641_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2584 <= data_out(223 downto 208);
      call1_2587 <= data_out(207 downto 192);
      call3_2590 <= data_out(191 downto 176);
      call5_2593 <= data_out(175 downto 160);
      call7_2596 <= data_out(159 downto 144);
      call9_2599 <= data_out(143 downto 128);
      call11_2602 <= data_out(127 downto 112);
      call13_2605 <= data_out(111 downto 96);
      call14_2608 <= data_out(95 downto 80);
      call15_2611 <= data_out(79 downto 64);
      call16_2624 <= data_out(63 downto 48);
      call18_2636 <= data_out(47 downto 32);
      call20_2639 <= data_out(31 downto 16);
      call22_2642 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2930_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2930_inst_req_0;
      WPIPE_Block3_done_2930_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2930_inst_req_1;
      WPIPE_Block3_done_2930_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2932_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_28_load_0_req_1 : boolean;
  signal LOAD_count_28_load_0_ack_1 : boolean;
  signal LOAD_count_28_load_0_req_0 : boolean;
  signal LOAD_count_28_load_0_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_29/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_sample_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_update_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/rr
      -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_0); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_sample_completed_
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/ra
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_ack
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_29/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_update_completed_
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_28_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_28_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_28_word_address_0 <= "0";
    -- equivalence LOAD_count_28_gather_scatter
    process(LOAD_count_28_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_28_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_28_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_28_load_0_req_0;
      LOAD_count_28_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_28_load_0_req_1;
      LOAD_count_28_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_28_word_address_0;
      LOAD_count_28_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
