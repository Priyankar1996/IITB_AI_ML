-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_36_load_0_req_0 : boolean;
  signal ptr_deref_36_load_0_ack_0 : boolean;
  signal ptr_deref_36_load_0_req_1 : boolean;
  signal ptr_deref_36_load_0_ack_1 : boolean;
  signal ptr_deref_48_load_0_req_0 : boolean;
  signal ptr_deref_48_load_0_ack_0 : boolean;
  signal ptr_deref_48_load_0_req_1 : boolean;
  signal ptr_deref_48_load_0_ack_1 : boolean;
  signal type_cast_172_inst_req_1 : boolean;
  signal type_cast_172_inst_ack_1 : boolean;
  signal type_cast_182_inst_req_0 : boolean;
  signal ptr_deref_60_load_0_req_0 : boolean;
  signal ptr_deref_60_load_0_ack_0 : boolean;
  signal ptr_deref_60_load_0_req_1 : boolean;
  signal ptr_deref_60_load_0_ack_1 : boolean;
  signal type_cast_74_inst_req_0 : boolean;
  signal type_cast_74_inst_ack_0 : boolean;
  signal type_cast_74_inst_req_1 : boolean;
  signal type_cast_74_inst_ack_1 : boolean;
  signal if_stmt_89_branch_req_0 : boolean;
  signal if_stmt_89_branch_ack_1 : boolean;
  signal if_stmt_89_branch_ack_0 : boolean;
  signal type_cast_108_inst_req_0 : boolean;
  signal type_cast_108_inst_ack_0 : boolean;
  signal type_cast_108_inst_req_1 : boolean;
  signal type_cast_108_inst_ack_1 : boolean;
  signal array_obj_ref_143_index_offset_req_0 : boolean;
  signal array_obj_ref_143_index_offset_ack_0 : boolean;
  signal array_obj_ref_143_index_offset_req_1 : boolean;
  signal array_obj_ref_143_index_offset_ack_1 : boolean;
  signal addr_of_144_final_reg_req_0 : boolean;
  signal addr_of_144_final_reg_ack_0 : boolean;
  signal addr_of_144_final_reg_req_1 : boolean;
  signal addr_of_144_final_reg_ack_1 : boolean;
  signal ptr_deref_148_load_0_req_0 : boolean;
  signal ptr_deref_148_load_0_ack_0 : boolean;
  signal ptr_deref_148_load_0_req_1 : boolean;
  signal ptr_deref_148_load_0_ack_1 : boolean;
  signal type_cast_152_inst_req_0 : boolean;
  signal type_cast_152_inst_ack_0 : boolean;
  signal type_cast_152_inst_req_1 : boolean;
  signal type_cast_152_inst_ack_1 : boolean;
  signal type_cast_162_inst_req_0 : boolean;
  signal type_cast_162_inst_ack_0 : boolean;
  signal type_cast_162_inst_req_1 : boolean;
  signal type_cast_162_inst_ack_1 : boolean;
  signal type_cast_172_inst_req_0 : boolean;
  signal type_cast_172_inst_ack_0 : boolean;
  signal type_cast_182_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_1 : boolean;
  signal type_cast_182_inst_ack_1 : boolean;
  signal type_cast_192_inst_req_0 : boolean;
  signal type_cast_192_inst_ack_0 : boolean;
  signal type_cast_192_inst_req_1 : boolean;
  signal type_cast_192_inst_ack_1 : boolean;
  signal type_cast_202_inst_req_0 : boolean;
  signal type_cast_202_inst_ack_0 : boolean;
  signal type_cast_202_inst_req_1 : boolean;
  signal type_cast_202_inst_ack_1 : boolean;
  signal type_cast_212_inst_req_0 : boolean;
  signal type_cast_212_inst_ack_0 : boolean;
  signal type_cast_212_inst_req_1 : boolean;
  signal type_cast_212_inst_ack_1 : boolean;
  signal type_cast_222_inst_req_0 : boolean;
  signal type_cast_222_inst_ack_0 : boolean;
  signal type_cast_222_inst_req_1 : boolean;
  signal type_cast_222_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_224_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_224_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_224_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_224_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_227_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_227_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_227_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_227_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_230_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_230_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_230_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_230_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_233_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_233_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_233_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_233_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_236_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_236_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_236_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_236_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_239_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_239_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_239_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_239_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_242_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_242_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_242_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_242_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_245_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_245_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_245_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_245_inst_ack_1 : boolean;
  signal if_stmt_259_branch_req_0 : boolean;
  signal if_stmt_259_branch_ack_1 : boolean;
  signal if_stmt_259_branch_ack_0 : boolean;
  signal phi_stmt_131_req_0 : boolean;
  signal type_cast_137_inst_req_0 : boolean;
  signal type_cast_137_inst_ack_0 : boolean;
  signal type_cast_137_inst_req_1 : boolean;
  signal type_cast_137_inst_ack_1 : boolean;
  signal phi_stmt_131_req_1 : boolean;
  signal phi_stmt_131_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(68);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (86) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_25/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/branch_block_stmt_25__entry__
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88__entry__
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_Update/cr
      -- 
    rr_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_36_load_0_req_0); -- 
    cr_100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_36_load_0_req_1); -- 
    rr_139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_48_load_0_req_0); -- 
    cr_150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_48_load_0_req_1); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_60_load_0_req_0); -- 
    cr_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_60_load_0_req_1); -- 
    cr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => type_cast_74_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Sample/word_access_start/word_0/ra
      -- 
    ra_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_36_load_0_ack_0, ack => sendOutput_CP_26_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/ptr_deref_36_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/ptr_deref_36_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/ptr_deref_36_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_36_Update/ptr_deref_36_Merge/merge_ack
      -- 
    ca_101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_36_load_0_ack_1, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Sample/word_access_start/word_0/ra
      -- 
    ra_140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_48_load_0_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/ptr_deref_48_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/ptr_deref_48_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/ptr_deref_48_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_48_Update/ptr_deref_48_Merge/merge_ack
      -- 
    ca_151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_48_load_0_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Sample/word_access_start/word_0/ra
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_60_load_0_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/ptr_deref_60_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/ptr_deref_60_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/ptr_deref_60_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/ptr_deref_60_Update/ptr_deref_60_Merge/merge_ack
      -- 
    ca_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_60_load_0_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_Sample/rr
      -- 
    rr_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(7), ack => type_cast_74_inst_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(2) & sendOutput_CP_26_elements(4) & sendOutput_CP_26_elements(6);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_Sample/ra
      -- 
    ra_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_74_inst_ack_0, ack => sendOutput_CP_26_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (13) 
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88__exit__
      -- CP-element group 9: 	 branch_block_stmt_25/if_stmt_89__entry__
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/$exit
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_33_to_assign_stmt_88/type_cast_74_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_25/if_stmt_89_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_25/if_stmt_89_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_25/if_stmt_89_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_25/if_stmt_89_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_25/R_cmp77_90_place
      -- CP-element group 9: 	 branch_block_stmt_25/if_stmt_89_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_25/if_stmt_89_else_link/$entry
      -- 
    ca_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_74_inst_ack_1, ack => sendOutput_CP_26_elements(9)); -- 
    branch_req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(9), ack => if_stmt_89_branch_req_0); -- 
    -- CP-element group 10:  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	68 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_25/if_stmt_89_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_25/if_stmt_89_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_25/entry_forx_xend
      -- CP-element group 10: 	 branch_block_stmt_25/entry_forx_xend_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_25/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_89_branch_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (18) 
      -- CP-element group 11: 	 branch_block_stmt_25/merge_stmt_95__exit__
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128__entry__
      -- CP-element group 11: 	 branch_block_stmt_25/if_stmt_89_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_25/if_stmt_89_else_link/else_choice_transition
      -- CP-element group 11: 	 branch_block_stmt_25/entry_bbx_xnph
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/$entry
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_update_start_
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_25/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_25/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_25/merge_stmt_95_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_25/merge_stmt_95_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_25/merge_stmt_95_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_25/merge_stmt_95_PhiAck/dummy
      -- 
    else_choice_transition_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_89_branch_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    rr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(11), ack => type_cast_108_inst_req_0); -- 
    cr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(11), ack => type_cast_108_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_Sample/ra
      -- 
    ra_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_108_inst_ack_0, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  place  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	62 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128__exit__
      -- CP-element group 13: 	 branch_block_stmt_25/bbx_xnph_forx_xbody
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/$exit
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_100_to_assign_stmt_128/type_cast_108_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_25/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_25/bbx_xnph_forx_xbody_PhiReq/phi_stmt_131/$entry
      -- CP-element group 13: 	 branch_block_stmt_25/bbx_xnph_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/$entry
      -- 
    ca_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_108_inst_ack_1, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	67 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	59 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_sample_complete
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_Sample/ack
      -- 
    ack_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_143_index_offset_ack_0, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	67 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (11) 
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_Update/ack
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_request/$entry
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_request/req
      -- 
    ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_143_index_offset_ack_1, ack => sendOutput_CP_26_elements(15)); -- 
    req_299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => addr_of_144_final_reg_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_request/$exit
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_request/ack
      -- 
    ack_300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_144_final_reg_ack_0, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	67 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (24) 
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_complete/ack
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_word_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_root_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_address_resized
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_addr_resize/$entry
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_addr_resize/$exit
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_addr_resize/base_resize_req
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_addr_resize/base_resize_ack
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_plus_offset/$entry
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_plus_offset/$exit
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_word_addrgen/$entry
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_word_addrgen/$exit
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_word_addrgen/root_register_req
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_word_addrgen/root_register_ack
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Sample/word_access_start/$entry
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Sample/word_access_start/word_0/$entry
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Sample/word_access_start/word_0/rr
      -- 
    ack_305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_144_final_reg_ack_1, ack => sendOutput_CP_26_elements(17)); -- 
    rr_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(17), ack => ptr_deref_148_load_0_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Sample/word_access_start/$exit
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Sample/word_access_start/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Sample/word_access_start/word_0/ra
      -- 
    ra_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_148_load_0_ack_0, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	67 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	26 
    -- CP-element group 19: 	28 
    -- CP-element group 19: 	30 
    -- CP-element group 19: 	32 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (33) 
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/word_access_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/word_access_complete/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/word_access_complete/word_0/ca
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/ptr_deref_148_Merge/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/ptr_deref_148_Merge/$exit
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/ptr_deref_148_Merge/merge_req
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/ptr_deref_148_Merge/merge_ack
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_Sample/rr
      -- 
    ca_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_148_load_0_ack_1, ack => sendOutput_CP_26_elements(19)); -- 
    rr_363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_152_inst_req_0); -- 
    rr_377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_162_inst_req_0); -- 
    rr_391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_172_inst_req_0); -- 
    rr_405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_182_inst_req_0); -- 
    rr_419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_192_inst_req_0); -- 
    rr_433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_202_inst_req_0); -- 
    rr_447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_212_inst_req_0); -- 
    rr_461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_222_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_Sample/ra
      -- 
    ra_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_0, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	67 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	56 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_Update/ca
      -- 
    ca_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_1, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_Sample/ra
      -- 
    ra_378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_162_inst_ack_0, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	67 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	53 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_Update/ca
      -- 
    ca_383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_162_inst_ack_1, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	19 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_Sample/ra
      -- 
    ra_392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_172_inst_ack_0, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	67 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_update_completed_
      -- 
    ca_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_172_inst_ack_1, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	19 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_Sample/ra
      -- 
    ra_406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_0, ack => sendOutput_CP_26_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	67 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	47 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_Update/ca
      -- 
    ca_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_1, ack => sendOutput_CP_26_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	19 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_Sample/ra
      -- 
    ra_420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_0, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	67 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	44 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_Update/ca
      -- 
    ca_425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_1, ack => sendOutput_CP_26_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	19 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_Sample/ra
      -- 
    ra_434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	67 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	41 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_Update/ca
      -- 
    ca_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	19 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_Sample/ra
      -- 
    ra_448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_0, ack => sendOutput_CP_26_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	67 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	38 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_Update/ca
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_1, ack => sendOutput_CP_26_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	19 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_Sample/ra
      -- 
    ra_462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_222_inst_ack_0, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	67 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_Sample/req
      -- 
    ca_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_222_inst_ack_1, ack => sendOutput_CP_26_elements(35)); -- 
    req_475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_224_inst_req_0); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_update_start_
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_Update/req
      -- 
    ack_476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_224_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_224_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_224_Update/ack
      -- 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_224_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	33 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_Sample/req
      -- 
    req_489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_227_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(33) & sendOutput_CP_26_elements(37);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_update_start_
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_Update/req
      -- 
    ack_490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_227_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_227_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_227_Update/ack
      -- 
    ack_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_227_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	31 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_Sample/req
      -- 
    req_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_230_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(31) & sendOutput_CP_26_elements(40);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_update_start_
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_Update/req
      -- 
    ack_504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_230_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_230_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_230_Update/ack
      -- 
    ack_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_230_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	29 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_Sample/req
      -- 
    req_517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_233_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(29) & sendOutput_CP_26_elements(43);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_update_start_
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_Update/req
      -- 
    ack_518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_233_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_233_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_233_Update/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_233_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	27 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_Sample/req
      -- 
    req_531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_236_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(27) & sendOutput_CP_26_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_update_start_
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_Update/req
      -- 
    ack_532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_236_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_236_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_236_Update/ack
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_236_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_Sample/req
      -- 
    req_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => WPIPE_zeropad_output_pipe_239_inst_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(25) & sendOutput_CP_26_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_update_start_
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_Update/req
      -- 
    ack_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_239_inst_ack_0, ack => sendOutput_CP_26_elements(51)); -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(51), ack => WPIPE_zeropad_output_pipe_239_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_239_Update/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_239_inst_ack_1, ack => sendOutput_CP_26_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	23 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_Sample/req
      -- 
    req_559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => WPIPE_zeropad_output_pipe_242_inst_req_0); -- 
    sendOutput_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(23) & sendOutput_CP_26_elements(52);
      gj_sendOutput_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_update_start_
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_Update/req
      -- 
    ack_560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_242_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(54), ack => WPIPE_zeropad_output_pipe_242_inst_req_1); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_242_Update/ack
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_242_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	21 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_Sample/req
      -- 
    req_573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => WPIPE_zeropad_output_pipe_245_inst_req_0); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(21) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_update_start_
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_Update/req
      -- 
    ack_574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_245_inst_ack_0, ack => sendOutput_CP_26_elements(57)); -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(57), ack => WPIPE_zeropad_output_pipe_245_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/WPIPE_zeropad_output_pipe_245_Update/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_245_inst_ack_1, ack => sendOutput_CP_26_elements(58)); -- 
    -- CP-element group 59:  branch  join  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	14 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (10) 
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258__exit__
      -- CP-element group 59: 	 branch_block_stmt_25/if_stmt_259__entry__
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/$exit
      -- CP-element group 59: 	 branch_block_stmt_25/if_stmt_259_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_25/if_stmt_259_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_25/if_stmt_259_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_25/if_stmt_259_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_25/R_exitcond9_260_place
      -- CP-element group 59: 	 branch_block_stmt_25/if_stmt_259_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_25/if_stmt_259_else_link/$entry
      -- 
    branch_req_587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(59), ack => if_stmt_259_branch_req_0); -- 
    sendOutput_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(14) & sendOutput_CP_26_elements(58);
      gj_sendOutput_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  merge  transition  place  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (13) 
      -- CP-element group 60: 	 branch_block_stmt_25/merge_stmt_265__exit__
      -- CP-element group 60: 	 branch_block_stmt_25/forx_xendx_xloopexit_forx_xend
      -- CP-element group 60: 	 branch_block_stmt_25/if_stmt_259_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_25/if_stmt_259_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_25/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 60: 	 branch_block_stmt_25/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_25/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_25/merge_stmt_265_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_25/merge_stmt_265_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_25/merge_stmt_265_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_25/merge_stmt_265_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_25/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_25/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_259_branch_ack_1, ack => sendOutput_CP_26_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	64 
    -- CP-element group 61:  members (12) 
      -- CP-element group 61: 	 branch_block_stmt_25/if_stmt_259_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_25/if_stmt_259_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/$entry
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/$entry
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/Update/cr
      -- 
    else_choice_transition_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_259_branch_ack_0, ack => sendOutput_CP_26_elements(61)); -- 
    rr_640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(61), ack => type_cast_137_inst_req_0); -- 
    cr_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(61), ack => type_cast_137_inst_req_1); -- 
    -- CP-element group 62:  transition  output  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	13 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	66 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_25/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_25/bbx_xnph_forx_xbody_PhiReq/phi_stmt_131/$exit
      -- CP-element group 62: 	 branch_block_stmt_25/bbx_xnph_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/$exit
      -- CP-element group 62: 	 branch_block_stmt_25/bbx_xnph_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_135_konst_delay_trans
      -- CP-element group 62: 	 branch_block_stmt_25/bbx_xnph_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_req
      -- 
    phi_stmt_131_req_621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_131_req_621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(62), ack => phi_stmt_131_req_0); -- 
    -- Element group sendOutput_CP_26_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(13), ack => sendOutput_CP_26_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/Sample/ra
      -- 
    ra_641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_137_inst_ack_0, ack => sendOutput_CP_26_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	61 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/Update/ca
      -- 
    ca_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_137_inst_ack_1, ack => sendOutput_CP_26_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/$exit
      -- CP-element group 65: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/$exit
      -- CP-element group 65: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_sources/type_cast_137/SplitProtocol/$exit
      -- CP-element group 65: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_131/phi_stmt_131_req
      -- 
    phi_stmt_131_req_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_131_req_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(65), ack => phi_stmt_131_req_1); -- 
    sendOutput_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(63) & sendOutput_CP_26_elements(64);
      gj_sendOutput_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_25/merge_stmt_130_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_25/merge_stmt_130_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(66) <= OrReduce(sendOutput_CP_26_elements(62) & sendOutput_CP_26_elements(65));
    -- CP-element group 67:  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: 	15 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	19 
    -- CP-element group 67: 	21 
    -- CP-element group 67: 	23 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	27 
    -- CP-element group 67: 	29 
    -- CP-element group 67: 	31 
    -- CP-element group 67: 	33 
    -- CP-element group 67: 	35 
    -- CP-element group 67:  members (53) 
      -- CP-element group 67: 	 branch_block_stmt_25/merge_stmt_130__exit__
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258__entry__
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_resized_1
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_scaled_1
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_computed_1
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_resize_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_resize_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_resize_1/index_resize_req
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_resize_1/index_resize_ack
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_scale_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_scale_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_scale_1/scale_rename_req
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_index_scale_1/scale_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_update_start
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/array_obj_ref_143_final_index_sum_regn_Update/req
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/addr_of_144_complete/req
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/word_access_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/word_access_complete/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/ptr_deref_148_Update/word_access_complete/word_0/cr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_152_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_162_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_172_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_182_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_192_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_202_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_212_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_update_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_145_to_assign_stmt_258/type_cast_222_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_25/merge_stmt_130_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_25/merge_stmt_130_PhiAck/phi_stmt_131_ack
      -- 
    phi_stmt_131_ack_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_131_ack_0, ack => sendOutput_CP_26_elements(67)); -- 
    cr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_172_inst_req_1); -- 
    req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => array_obj_ref_143_index_offset_req_0); -- 
    req_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => array_obj_ref_143_index_offset_req_1); -- 
    req_304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => addr_of_144_final_reg_req_1); -- 
    cr_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => ptr_deref_148_load_0_req_1); -- 
    cr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_152_inst_req_1); -- 
    cr_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_162_inst_req_1); -- 
    cr_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_182_inst_req_1); -- 
    cr_424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_192_inst_req_1); -- 
    cr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_202_inst_req_1); -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_212_inst_req_1); -- 
    cr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_222_inst_req_1); -- 
    -- CP-element group 68:  merge  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	10 
    -- CP-element group 68: 	60 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_25/$exit
      -- CP-element group 68: 	 branch_block_stmt_25/branch_block_stmt_25__exit__
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_267__exit__
      -- CP-element group 68: 	 branch_block_stmt_25/return__
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_269__exit__
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_267_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_267_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_267_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_267_PhiAck/dummy
      -- CP-element group 68: 	 branch_block_stmt_25/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_25/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_269_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_269_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_269_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_25/merge_stmt_269_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(68) <= OrReduce(sendOutput_CP_26_elements(10) & sendOutput_CP_26_elements(60));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_142_resized : std_logic_vector(13 downto 0);
    signal R_indvar_142_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_143_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_143_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_143_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_143_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_143_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_143_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_145 : std_logic_vector(31 downto 0);
    signal cmp77_88 : std_logic_vector(0 downto 0);
    signal conv14_153 : std_logic_vector(7 downto 0);
    signal conv20_163 : std_logic_vector(7 downto 0);
    signal conv26_173 : std_logic_vector(7 downto 0);
    signal conv32_183 : std_logic_vector(7 downto 0);
    signal conv38_193 : std_logic_vector(7 downto 0);
    signal conv44_203 : std_logic_vector(7 downto 0);
    signal conv50_213 : std_logic_vector(7 downto 0);
    signal conv56_223 : std_logic_vector(7 downto 0);
    signal conv_75 : std_logic_vector(63 downto 0);
    signal exitcond9_258 : std_logic_vector(0 downto 0);
    signal iNsTr_0_33 : std_logic_vector(31 downto 0);
    signal iNsTr_1_45 : std_logic_vector(31 downto 0);
    signal iNsTr_2_57 : std_logic_vector(31 downto 0);
    signal indvar_131 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_253 : std_logic_vector(63 downto 0);
    signal mul3_71 : std_logic_vector(31 downto 0);
    signal mul_66 : std_logic_vector(31 downto 0);
    signal ptr_deref_148_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_148_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_148_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_148_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_148_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_36_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_36_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_36_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_36_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_36_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_48_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_48_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_48_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_48_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_48_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_60_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_60_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_60_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_60_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_60_word_offset_0 : std_logic_vector(6 downto 0);
    signal shr17_159 : std_logic_vector(63 downto 0);
    signal shr23_169 : std_logic_vector(63 downto 0);
    signal shr29_179 : std_logic_vector(63 downto 0);
    signal shr35_189 : std_logic_vector(63 downto 0);
    signal shr41_199 : std_logic_vector(63 downto 0);
    signal shr47_209 : std_logic_vector(63 downto 0);
    signal shr53_219 : std_logic_vector(63 downto 0);
    signal shr76x_xmask_81 : std_logic_vector(63 downto 0);
    signal tmp11_149 : std_logic_vector(63 downto 0);
    signal tmp1_49 : std_logic_vector(31 downto 0);
    signal tmp2_61 : std_logic_vector(31 downto 0);
    signal tmp3_100 : std_logic_vector(31 downto 0);
    signal tmp4_105 : std_logic_vector(31 downto 0);
    signal tmp5_109 : std_logic_vector(63 downto 0);
    signal tmp6_115 : std_logic_vector(63 downto 0);
    signal tmp7_121 : std_logic_vector(0 downto 0);
    signal tmp_37 : std_logic_vector(31 downto 0);
    signal type_cast_113_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_119_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_126_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_135_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_137_wire : std_logic_vector(63 downto 0);
    signal type_cast_157_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_167_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_177_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_187_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_197_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_207_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_217_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_251_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_79_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_85_wire_constant : std_logic_vector(63 downto 0);
    signal umax8_128 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_143_constant_part_of_offset <= "00000000000000";
    array_obj_ref_143_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_143_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_143_resized_base_address <= "00000000000000";
    iNsTr_0_33 <= "00000000000000000000000000000010";
    iNsTr_1_45 <= "00000000000000000000000000000011";
    iNsTr_2_57 <= "00000000000000000000000000000100";
    ptr_deref_148_word_offset_0 <= "00000000000000";
    ptr_deref_36_word_offset_0 <= "0000000";
    ptr_deref_48_word_offset_0 <= "0000000";
    ptr_deref_60_word_offset_0 <= "0000000";
    type_cast_113_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_119_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_126_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_135_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_157_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_167_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_177_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_187_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_197_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_207_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_217_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_251_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_79_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_85_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_131: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_135_wire_constant & type_cast_137_wire;
      req <= phi_stmt_131_req_0 & phi_stmt_131_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_131",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_131_ack_0,
          idata => idata,
          odata => indvar_131,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_131
    -- flow-through select operator MUX_127_inst
    umax8_128 <= tmp6_115 when (tmp7_121(0) /=  '0') else type_cast_126_wire_constant;
    addr_of_144_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_144_final_reg_req_0;
      addr_of_144_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_144_final_reg_req_1;
      addr_of_144_final_reg_ack_1<= rack(0);
      addr_of_144_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_144_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_143_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_108_inst_req_0;
      type_cast_108_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_108_inst_req_1;
      type_cast_108_inst_ack_1<= rack(0);
      type_cast_108_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_105,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp5_109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_137_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_137_inst_req_0;
      type_cast_137_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_137_inst_req_1;
      type_cast_137_inst_ack_1<= rack(0);
      type_cast_137_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_137_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_137_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_152_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_152_inst_req_0;
      type_cast_152_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_152_inst_req_1;
      type_cast_152_inst_ack_1<= rack(0);
      type_cast_152_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_152_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_162_inst_req_0;
      type_cast_162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_162_inst_req_1;
      type_cast_162_inst_ack_1<= rack(0);
      type_cast_162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_159,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_163,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_172_inst_req_0;
      type_cast_172_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_172_inst_req_1;
      type_cast_172_inst_ack_1<= rack(0);
      type_cast_172_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_172_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_169,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_182_inst_req_0;
      type_cast_182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_182_inst_req_1;
      type_cast_182_inst_ack_1<= rack(0);
      type_cast_182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_192_inst_req_0;
      type_cast_192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_192_inst_req_1;
      type_cast_192_inst_ack_1<= rack(0);
      type_cast_192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_202_inst_req_0;
      type_cast_202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_202_inst_req_1;
      type_cast_202_inst_ack_1<= rack(0);
      type_cast_202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_212_inst_req_0;
      type_cast_212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_212_inst_req_1;
      type_cast_212_inst_ack_1<= rack(0);
      type_cast_212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr47_209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_222_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_222_inst_req_0;
      type_cast_222_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_222_inst_req_1;
      type_cast_222_inst_ack_1<= rack(0);
      type_cast_222_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_222_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr53_219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_74_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_74_inst_req_0;
      type_cast_74_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_74_inst_req_1;
      type_cast_74_inst_ack_1<= rack(0);
      type_cast_74_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_74_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul3_71,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_75,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_143_index_1_rename
    process(R_indvar_142_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_142_resized;
      ov(13 downto 0) := iv;
      R_indvar_142_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_143_index_1_resize
    process(indvar_131) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_131;
      ov := iv(13 downto 0);
      R_indvar_142_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_143_root_address_inst
    process(array_obj_ref_143_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_143_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_143_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_148_addr_0
    process(ptr_deref_148_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_148_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_148_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_148_base_resize
    process(arrayidx_145) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_145;
      ov := iv(13 downto 0);
      ptr_deref_148_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_148_gather_scatter
    process(ptr_deref_148_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_148_data_0;
      ov(63 downto 0) := iv;
      tmp11_149 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_148_root_address_inst
    process(ptr_deref_148_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_148_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_148_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_36_addr_0
    process(ptr_deref_36_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_36_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_36_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_36_base_resize
    process(iNsTr_0_33) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_33;
      ov := iv(6 downto 0);
      ptr_deref_36_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_36_gather_scatter
    process(ptr_deref_36_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_36_data_0;
      ov(31 downto 0) := iv;
      tmp_37 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_36_root_address_inst
    process(ptr_deref_36_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_36_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_36_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_48_addr_0
    process(ptr_deref_48_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_48_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_48_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_48_base_resize
    process(iNsTr_1_45) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_45;
      ov := iv(6 downto 0);
      ptr_deref_48_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_48_gather_scatter
    process(ptr_deref_48_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_48_data_0;
      ov(31 downto 0) := iv;
      tmp1_49 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_48_root_address_inst
    process(ptr_deref_48_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_48_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_48_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_60_addr_0
    process(ptr_deref_60_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_60_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_60_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_60_base_resize
    process(iNsTr_2_57) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_57;
      ov := iv(6 downto 0);
      ptr_deref_60_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_60_gather_scatter
    process(ptr_deref_60_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_60_data_0;
      ov(31 downto 0) := iv;
      tmp2_61 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_60_root_address_inst
    process(ptr_deref_60_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_60_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_60_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_259_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond9_258;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_259_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_259_branch_req_0,
          ack0 => if_stmt_259_branch_ack_0,
          ack1 => if_stmt_259_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_89_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_88;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_89_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_89_branch_req_0,
          ack0 => if_stmt_89_branch_ack_0,
          ack1 => if_stmt_89_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_252_inst
    process(indvar_131) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_131, type_cast_251_wire_constant, tmp_var);
      indvarx_xnext_253 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_80_inst
    process(conv_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv_75, type_cast_79_wire_constant, tmp_var);
      shr76x_xmask_81 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_257_inst
    process(indvarx_xnext_253, umax8_128) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_253, umax8_128, tmp_var);
      exitcond9_258 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_86_inst
    process(shr76x_xmask_81) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr76x_xmask_81, type_cast_85_wire_constant, tmp_var);
      cmp77_88 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_114_inst
    process(tmp5_109) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_109, type_cast_113_wire_constant, tmp_var);
      tmp6_115 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_158_inst
    process(tmp11_149) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_149, type_cast_157_wire_constant, tmp_var);
      shr17_159 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_168_inst
    process(tmp11_149) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_149, type_cast_167_wire_constant, tmp_var);
      shr23_169 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_178_inst
    process(tmp11_149) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_149, type_cast_177_wire_constant, tmp_var);
      shr29_179 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_188_inst
    process(tmp11_149) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_149, type_cast_187_wire_constant, tmp_var);
      shr35_189 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_198_inst
    process(tmp11_149) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_149, type_cast_197_wire_constant, tmp_var);
      shr41_199 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_208_inst
    process(tmp11_149) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_149, type_cast_207_wire_constant, tmp_var);
      shr47_209 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_218_inst
    process(tmp11_149) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_149, type_cast_217_wire_constant, tmp_var);
      shr53_219 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_104_inst
    process(tmp3_100, tmp2_61) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_100, tmp2_61, tmp_var);
      tmp4_105 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_65_inst
    process(tmp1_49, tmp_37) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_49, tmp_37, tmp_var);
      mul_66 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_70_inst
    process(mul_66, tmp2_61) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_66, tmp2_61, tmp_var);
      mul3_71 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_99_inst
    process(tmp1_49, tmp_37) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_49, tmp_37, tmp_var);
      tmp3_100 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_120_inst
    process(tmp6_115) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp6_115, type_cast_119_wire_constant, tmp_var);
      tmp7_121 <= tmp_var; --
    end process;
    -- shared split operator group (17) : array_obj_ref_143_index_offset 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_142_scaled;
      array_obj_ref_143_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_143_index_offset_req_0;
      array_obj_ref_143_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_143_index_offset_req_1;
      array_obj_ref_143_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared load operator group (0) : ptr_deref_148_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_148_load_0_req_0;
      ptr_deref_148_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_148_load_0_req_1;
      ptr_deref_148_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_148_word_address_0;
      ptr_deref_148_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_36_load_0 ptr_deref_48_load_0 ptr_deref_60_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_36_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_48_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_60_load_0_req_0;
      ptr_deref_36_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_48_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_60_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_36_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_48_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_60_load_0_req_1;
      ptr_deref_36_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_48_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_60_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_36_word_address_0 & ptr_deref_48_word_address_0 & ptr_deref_60_word_address_0;
      ptr_deref_36_data_0 <= data_out(95 downto 64);
      ptr_deref_48_data_0 <= data_out(63 downto 32);
      ptr_deref_60_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_224_inst WPIPE_zeropad_output_pipe_227_inst WPIPE_zeropad_output_pipe_230_inst WPIPE_zeropad_output_pipe_233_inst WPIPE_zeropad_output_pipe_236_inst WPIPE_zeropad_output_pipe_239_inst WPIPE_zeropad_output_pipe_242_inst WPIPE_zeropad_output_pipe_245_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_224_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_227_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_230_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_233_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_236_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_239_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_242_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_245_inst_req_0;
      WPIPE_zeropad_output_pipe_224_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_227_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_230_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_233_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_236_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_239_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_242_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_245_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_224_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_227_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_230_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_233_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_236_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_239_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_242_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_245_inst_req_1;
      WPIPE_zeropad_output_pipe_224_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_227_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_230_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_233_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_236_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_239_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_242_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_245_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv56_223 & conv50_213 & conv44_203 & conv38_193 & conv32_183 & conv26_173 & conv20_163 & conv14_153;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(8 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_684_start: Boolean;
  signal testConfigure_CP_684_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_314_addr_3_req_1 : boolean;
  signal ptr_deref_489_addr_3_ack_1 : boolean;
  signal ptr_deref_314_addr_3_req_0 : boolean;
  signal ptr_deref_501_addr_3_ack_1 : boolean;
  signal ptr_deref_314_addr_3_ack_1 : boolean;
  signal ptr_deref_314_addr_3_ack_0 : boolean;
  signal ptr_deref_314_addr_2_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_301_inst_ack_1 : boolean;
  signal type_cast_305_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_288_inst_ack_1 : boolean;
  signal ptr_deref_489_load_0_req_0 : boolean;
  signal ptr_deref_283_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_288_inst_ack_0 : boolean;
  signal ptr_deref_283_addr_3_ack_0 : boolean;
  signal ptr_deref_489_load_3_req_0 : boolean;
  signal ptr_deref_297_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_301_inst_req_1 : boolean;
  signal ptr_deref_297_store_0_req_1 : boolean;
  signal ptr_deref_314_addr_1_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_288_inst_req_0 : boolean;
  signal ptr_deref_314_addr_1_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_288_inst_req_1 : boolean;
  signal type_cast_305_inst_req_1 : boolean;
  signal ptr_deref_283_addr_3_req_0 : boolean;
  signal ptr_deref_501_load_2_req_0 : boolean;
  signal ptr_deref_489_load_2_req_0 : boolean;
  signal ptr_deref_314_addr_1_req_1 : boolean;
  signal ptr_deref_489_load_2_ack_0 : boolean;
  signal ptr_deref_314_addr_0_ack_1 : boolean;
  signal ptr_deref_283_addr_2_ack_1 : boolean;
  signal ptr_deref_283_addr_2_req_1 : boolean;
  signal ptr_deref_314_addr_0_req_1 : boolean;
  signal ptr_deref_297_store_0_req_0 : boolean;
  signal ptr_deref_283_store_3_ack_1 : boolean;
  signal ptr_deref_283_store_3_req_1 : boolean;
  signal ptr_deref_283_addr_2_ack_0 : boolean;
  signal type_cast_305_inst_ack_0 : boolean;
  signal ptr_deref_283_addr_2_req_0 : boolean;
  signal ptr_deref_314_addr_2_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_301_inst_ack_0 : boolean;
  signal ptr_deref_457_store_0_req_0 : boolean;
  signal type_cast_305_inst_req_0 : boolean;
  signal ptr_deref_283_store_2_ack_1 : boolean;
  signal ptr_deref_457_store_0_ack_0 : boolean;
  signal ptr_deref_283_addr_1_ack_1 : boolean;
  signal ptr_deref_283_addr_1_req_1 : boolean;
  signal ptr_deref_283_store_2_req_1 : boolean;
  signal ptr_deref_489_load_3_ack_0 : boolean;
  signal ptr_deref_283_store_1_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_301_inst_req_0 : boolean;
  signal ptr_deref_314_addr_0_ack_0 : boolean;
  signal ptr_deref_489_load_0_ack_0 : boolean;
  signal ptr_deref_314_addr_0_req_0 : boolean;
  signal ptr_deref_489_load_1_ack_0 : boolean;
  signal ptr_deref_283_addr_1_ack_0 : boolean;
  signal ptr_deref_283_addr_1_req_0 : boolean;
  signal ptr_deref_283_store_1_req_1 : boolean;
  signal ptr_deref_501_load_2_ack_0 : boolean;
  signal ptr_deref_283_store_0_ack_1 : boolean;
  signal ptr_deref_283_store_0_req_1 : boolean;
  signal ptr_deref_283_addr_3_ack_1 : boolean;
  signal ptr_deref_283_addr_0_ack_1 : boolean;
  signal ptr_deref_283_addr_0_req_1 : boolean;
  signal ptr_deref_283_addr_0_ack_0 : boolean;
  signal ptr_deref_283_addr_0_req_0 : boolean;
  signal ptr_deref_297_store_0_ack_0 : boolean;
  signal ptr_deref_283_store_3_ack_0 : boolean;
  signal ptr_deref_283_store_3_req_0 : boolean;
  signal ptr_deref_513_addr_2_req_1 : boolean;
  signal ptr_deref_513_addr_1_ack_0 : boolean;
  signal ptr_deref_513_load_0_req_0 : boolean;
  signal ptr_deref_501_load_3_req_1 : boolean;
  signal ptr_deref_501_load_3_ack_1 : boolean;
  signal ptr_deref_513_addr_2_ack_1 : boolean;
  signal ptr_deref_283_store_2_ack_0 : boolean;
  signal ptr_deref_283_store_2_req_0 : boolean;
  signal ptr_deref_283_store_1_ack_0 : boolean;
  signal ptr_deref_283_store_1_req_0 : boolean;
  signal ptr_deref_489_load_1_req_0 : boolean;
  signal ptr_deref_501_load_1_req_1 : boolean;
  signal ptr_deref_314_addr_2_ack_0 : boolean;
  signal ptr_deref_314_addr_2_req_0 : boolean;
  signal ptr_deref_314_addr_1_ack_0 : boolean;
  signal ptr_deref_283_store_0_ack_0 : boolean;
  signal ptr_deref_501_load_3_req_0 : boolean;
  signal ptr_deref_476_store_0_req_1 : boolean;
  signal ptr_deref_476_store_0_ack_1 : boolean;
  signal ptr_deref_489_load_0_req_1 : boolean;
  signal ptr_deref_501_load_2_req_1 : boolean;
  signal ptr_deref_501_load_3_ack_0 : boolean;
  signal ptr_deref_489_load_0_ack_1 : boolean;
  signal ptr_deref_501_load_0_req_0 : boolean;
  signal ptr_deref_457_store_0_req_1 : boolean;
  signal ptr_deref_513_addr_0_req_0 : boolean;
  signal ptr_deref_513_load_0_ack_0 : boolean;
  signal ptr_deref_513_load_3_req_0 : boolean;
  signal ptr_deref_501_load_2_ack_1 : boolean;
  signal ptr_deref_513_addr_3_req_1 : boolean;
  signal ptr_deref_513_load_1_req_0 : boolean;
  signal ptr_deref_513_load_0_req_1 : boolean;
  signal ptr_deref_513_load_0_ack_1 : boolean;
  signal ptr_deref_513_load_1_ack_0 : boolean;
  signal ptr_deref_513_load_2_req_0 : boolean;
  signal ptr_deref_513_load_2_ack_0 : boolean;
  signal ptr_deref_513_addr_1_req_0 : boolean;
  signal ptr_deref_513_addr_3_ack_1 : boolean;
  signal ptr_deref_513_addr_2_req_0 : boolean;
  signal ptr_deref_513_addr_2_ack_0 : boolean;
  signal ptr_deref_513_addr_0_ack_0 : boolean;
  signal ptr_deref_513_addr_3_req_0 : boolean;
  signal ptr_deref_513_addr_3_ack_0 : boolean;
  signal ptr_deref_513_addr_1_req_1 : boolean;
  signal ptr_deref_513_load_3_ack_0 : boolean;
  signal ptr_deref_457_store_0_ack_1 : boolean;
  signal ptr_deref_489_load_1_req_1 : boolean;
  signal ptr_deref_489_load_1_ack_1 : boolean;
  signal ptr_deref_501_load_1_ack_1 : boolean;
  signal ptr_deref_513_addr_1_ack_1 : boolean;
  signal ptr_deref_476_store_0_req_0 : boolean;
  signal ptr_deref_489_load_2_req_1 : boolean;
  signal ptr_deref_513_addr_0_req_1 : boolean;
  signal ptr_deref_489_load_2_ack_1 : boolean;
  signal ptr_deref_476_store_0_ack_0 : boolean;
  signal ptr_deref_489_load_3_req_1 : boolean;
  signal ptr_deref_489_load_3_ack_1 : boolean;
  signal ptr_deref_283_addr_3_req_1 : boolean;
  signal ptr_deref_314_store_0_req_0 : boolean;
  signal ptr_deref_314_store_0_ack_0 : boolean;
  signal ptr_deref_501_addr_3_req_1 : boolean;
  signal ptr_deref_314_store_1_req_0 : boolean;
  signal ptr_deref_314_store_1_ack_0 : boolean;
  signal ptr_deref_314_store_2_req_0 : boolean;
  signal ptr_deref_314_store_2_ack_0 : boolean;
  signal ptr_deref_314_store_3_req_0 : boolean;
  signal ptr_deref_314_store_3_ack_0 : boolean;
  signal ptr_deref_314_store_0_req_1 : boolean;
  signal ptr_deref_501_addr_3_ack_0 : boolean;
  signal ptr_deref_314_store_0_ack_1 : boolean;
  signal ptr_deref_489_addr_3_req_1 : boolean;
  signal ptr_deref_314_store_1_req_1 : boolean;
  signal ptr_deref_501_addr_3_req_0 : boolean;
  signal ptr_deref_314_store_1_ack_1 : boolean;
  signal ptr_deref_314_store_2_req_1 : boolean;
  signal ptr_deref_314_store_2_ack_1 : boolean;
  signal ptr_deref_314_store_3_req_1 : boolean;
  signal ptr_deref_314_store_3_ack_1 : boolean;
  signal ptr_deref_501_addr_2_ack_1 : boolean;
  signal ptr_deref_501_load_1_ack_0 : boolean;
  signal ptr_deref_501_load_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_req_0 : boolean;
  signal ptr_deref_501_addr_2_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_ack_1 : boolean;
  signal ptr_deref_489_addr_3_ack_0 : boolean;
  signal ptr_deref_489_addr_3_req_0 : boolean;
  signal ptr_deref_513_addr_0_ack_1 : boolean;
  signal ptr_deref_501_load_0_req_1 : boolean;
  signal type_cast_465_inst_ack_1 : boolean;
  signal if_stmt_326_branch_req_0 : boolean;
  signal ptr_deref_489_addr_2_ack_1 : boolean;
  signal if_stmt_326_branch_ack_1 : boolean;
  signal if_stmt_326_branch_ack_0 : boolean;
  signal ptr_deref_489_addr_2_req_1 : boolean;
  signal type_cast_357_inst_req_0 : boolean;
  signal ptr_deref_501_addr_2_ack_0 : boolean;
  signal type_cast_357_inst_ack_0 : boolean;
  signal type_cast_357_inst_req_1 : boolean;
  signal ptr_deref_501_addr_2_req_0 : boolean;
  signal type_cast_357_inst_ack_1 : boolean;
  signal type_cast_465_inst_req_1 : boolean;
  signal ptr_deref_501_load_1_req_0 : boolean;
  signal ptr_deref_489_addr_2_ack_0 : boolean;
  signal ptr_deref_489_addr_2_req_0 : boolean;
  signal ptr_deref_489_addr_1_ack_1 : boolean;
  signal ptr_deref_489_addr_1_req_1 : boolean;
  signal array_obj_ref_363_index_1_scale_req_0 : boolean;
  signal array_obj_ref_363_index_1_scale_ack_0 : boolean;
  signal array_obj_ref_363_index_1_scale_req_1 : boolean;
  signal array_obj_ref_363_index_1_scale_ack_1 : boolean;
  signal type_cast_465_inst_ack_0 : boolean;
  signal array_obj_ref_363_index_offset_req_0 : boolean;
  signal array_obj_ref_363_index_offset_ack_0 : boolean;
  signal type_cast_465_inst_req_0 : boolean;
  signal array_obj_ref_363_index_offset_req_1 : boolean;
  signal ptr_deref_501_addr_1_ack_1 : boolean;
  signal array_obj_ref_363_index_offset_ack_1 : boolean;
  signal ptr_deref_501_addr_1_req_1 : boolean;
  signal addr_of_364_final_reg_req_0 : boolean;
  signal addr_of_364_final_reg_ack_0 : boolean;
  signal addr_of_364_final_reg_req_1 : boolean;
  signal ptr_deref_501_addr_1_ack_0 : boolean;
  signal addr_of_364_final_reg_ack_1 : boolean;
  signal ptr_deref_489_addr_1_ack_0 : boolean;
  signal ptr_deref_489_addr_1_req_0 : boolean;
  signal type_cast_368_inst_req_0 : boolean;
  signal ptr_deref_501_addr_1_req_0 : boolean;
  signal type_cast_368_inst_ack_0 : boolean;
  signal type_cast_368_inst_req_1 : boolean;
  signal type_cast_368_inst_ack_1 : boolean;
  signal ptr_deref_501_load_0_ack_0 : boolean;
  signal ptr_deref_489_addr_0_ack_1 : boolean;
  signal ptr_deref_489_addr_0_req_1 : boolean;
  signal ptr_deref_489_addr_0_ack_0 : boolean;
  signal ptr_deref_489_addr_0_req_0 : boolean;
  signal ptr_deref_501_addr_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_461_inst_ack_1 : boolean;
  signal ptr_deref_371_addr_0_req_0 : boolean;
  signal ptr_deref_501_addr_0_req_1 : boolean;
  signal ptr_deref_371_addr_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_461_inst_req_1 : boolean;
  signal ptr_deref_371_addr_0_req_1 : boolean;
  signal ptr_deref_371_addr_0_ack_1 : boolean;
  signal ptr_deref_371_addr_1_req_0 : boolean;
  signal ptr_deref_371_addr_1_ack_0 : boolean;
  signal ptr_deref_371_addr_1_req_1 : boolean;
  signal ptr_deref_501_addr_0_ack_0 : boolean;
  signal ptr_deref_371_addr_1_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_461_inst_ack_0 : boolean;
  signal ptr_deref_371_addr_2_req_0 : boolean;
  signal ptr_deref_501_addr_0_req_0 : boolean;
  signal ptr_deref_371_addr_2_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_461_inst_req_0 : boolean;
  signal ptr_deref_371_addr_2_req_1 : boolean;
  signal ptr_deref_371_addr_2_ack_1 : boolean;
  signal ptr_deref_371_addr_3_req_0 : boolean;
  signal ptr_deref_371_addr_3_ack_0 : boolean;
  signal ptr_deref_371_addr_3_req_1 : boolean;
  signal ptr_deref_371_addr_3_ack_1 : boolean;
  signal ptr_deref_371_store_0_req_0 : boolean;
  signal ptr_deref_371_store_0_ack_0 : boolean;
  signal ptr_deref_371_store_1_req_0 : boolean;
  signal ptr_deref_371_store_1_ack_0 : boolean;
  signal ptr_deref_371_store_2_req_0 : boolean;
  signal ptr_deref_371_store_2_ack_0 : boolean;
  signal ptr_deref_371_store_3_req_0 : boolean;
  signal ptr_deref_371_store_3_ack_0 : boolean;
  signal ptr_deref_371_store_0_req_1 : boolean;
  signal ptr_deref_371_store_0_ack_1 : boolean;
  signal ptr_deref_371_store_1_req_1 : boolean;
  signal ptr_deref_371_store_1_ack_1 : boolean;
  signal ptr_deref_371_store_2_req_1 : boolean;
  signal ptr_deref_371_store_2_ack_1 : boolean;
  signal ptr_deref_371_store_3_req_1 : boolean;
  signal ptr_deref_371_store_3_ack_1 : boolean;
  signal ptr_deref_388_addr_0_req_0 : boolean;
  signal ptr_deref_388_addr_0_ack_0 : boolean;
  signal ptr_deref_388_addr_0_req_1 : boolean;
  signal ptr_deref_388_addr_0_ack_1 : boolean;
  signal ptr_deref_388_addr_1_req_0 : boolean;
  signal ptr_deref_388_addr_1_ack_0 : boolean;
  signal ptr_deref_388_addr_1_req_1 : boolean;
  signal ptr_deref_388_addr_1_ack_1 : boolean;
  signal ptr_deref_388_addr_2_req_0 : boolean;
  signal ptr_deref_388_addr_2_ack_0 : boolean;
  signal ptr_deref_388_addr_2_req_1 : boolean;
  signal ptr_deref_388_addr_2_ack_1 : boolean;
  signal ptr_deref_388_addr_3_req_0 : boolean;
  signal ptr_deref_388_addr_3_ack_0 : boolean;
  signal ptr_deref_388_addr_3_req_1 : boolean;
  signal ptr_deref_388_addr_3_ack_1 : boolean;
  signal ptr_deref_388_load_0_req_0 : boolean;
  signal ptr_deref_388_load_0_ack_0 : boolean;
  signal ptr_deref_388_load_1_req_0 : boolean;
  signal ptr_deref_388_load_1_ack_0 : boolean;
  signal ptr_deref_388_load_2_req_0 : boolean;
  signal ptr_deref_388_load_2_ack_0 : boolean;
  signal ptr_deref_388_load_3_req_0 : boolean;
  signal ptr_deref_388_load_3_ack_0 : boolean;
  signal ptr_deref_388_load_0_req_1 : boolean;
  signal ptr_deref_388_load_0_ack_1 : boolean;
  signal ptr_deref_388_load_1_req_1 : boolean;
  signal ptr_deref_388_load_1_ack_1 : boolean;
  signal ptr_deref_388_load_2_req_1 : boolean;
  signal ptr_deref_388_load_2_ack_1 : boolean;
  signal ptr_deref_388_load_3_req_1 : boolean;
  signal ptr_deref_388_load_3_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_396_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_396_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_396_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_396_inst_ack_1 : boolean;
  signal if_stmt_398_branch_req_0 : boolean;
  signal if_stmt_398_branch_ack_1 : boolean;
  signal if_stmt_398_branch_ack_0 : boolean;
  signal STORE_pad_419_store_0_req_0 : boolean;
  signal STORE_pad_419_store_0_ack_0 : boolean;
  signal STORE_pad_419_store_0_req_1 : boolean;
  signal STORE_pad_419_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_423_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_423_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_423_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_423_inst_ack_1 : boolean;
  signal type_cast_427_inst_req_0 : boolean;
  signal type_cast_427_inst_ack_0 : boolean;
  signal type_cast_427_inst_req_1 : boolean;
  signal type_cast_427_inst_ack_1 : boolean;
  signal ptr_deref_438_store_0_req_0 : boolean;
  signal ptr_deref_438_store_0_ack_0 : boolean;
  signal ptr_deref_438_store_0_req_1 : boolean;
  signal ptr_deref_438_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_442_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_442_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_442_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_442_inst_ack_1 : boolean;
  signal type_cast_446_inst_req_0 : boolean;
  signal type_cast_446_inst_ack_0 : boolean;
  signal type_cast_446_inst_req_1 : boolean;
  signal type_cast_446_inst_ack_1 : boolean;
  signal ptr_deref_513_load_1_req_1 : boolean;
  signal ptr_deref_513_load_1_ack_1 : boolean;
  signal ptr_deref_513_load_2_req_1 : boolean;
  signal ptr_deref_513_load_2_ack_1 : boolean;
  signal ptr_deref_513_load_3_req_1 : boolean;
  signal ptr_deref_513_load_3_ack_1 : boolean;
  signal type_cast_527_inst_req_0 : boolean;
  signal type_cast_527_inst_ack_0 : boolean;
  signal type_cast_527_inst_req_1 : boolean;
  signal type_cast_527_inst_ack_1 : boolean;
  signal if_stmt_541_branch_req_0 : boolean;
  signal if_stmt_541_branch_ack_1 : boolean;
  signal if_stmt_541_branch_ack_0 : boolean;
  signal type_cast_560_inst_req_0 : boolean;
  signal type_cast_560_inst_ack_0 : boolean;
  signal type_cast_560_inst_req_1 : boolean;
  signal type_cast_560_inst_ack_1 : boolean;
  signal array_obj_ref_595_index_offset_req_0 : boolean;
  signal array_obj_ref_595_index_offset_ack_0 : boolean;
  signal array_obj_ref_595_index_offset_req_1 : boolean;
  signal array_obj_ref_595_index_offset_ack_1 : boolean;
  signal addr_of_596_final_reg_req_0 : boolean;
  signal addr_of_596_final_reg_ack_0 : boolean;
  signal addr_of_596_final_reg_req_1 : boolean;
  signal addr_of_596_final_reg_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_599_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_599_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_599_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_599_inst_ack_1 : boolean;
  signal type_cast_603_inst_req_0 : boolean;
  signal type_cast_603_inst_ack_0 : boolean;
  signal type_cast_603_inst_req_1 : boolean;
  signal type_cast_603_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_612_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_612_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_612_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_612_inst_ack_1 : boolean;
  signal type_cast_616_inst_req_0 : boolean;
  signal type_cast_616_inst_ack_0 : boolean;
  signal type_cast_616_inst_req_1 : boolean;
  signal type_cast_616_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_630_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_630_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_630_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_630_inst_ack_1 : boolean;
  signal type_cast_634_inst_req_0 : boolean;
  signal type_cast_634_inst_ack_0 : boolean;
  signal type_cast_634_inst_req_1 : boolean;
  signal type_cast_634_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_648_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_648_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_648_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_648_inst_ack_1 : boolean;
  signal type_cast_652_inst_req_0 : boolean;
  signal type_cast_652_inst_ack_0 : boolean;
  signal type_cast_652_inst_req_1 : boolean;
  signal type_cast_652_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_666_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_666_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_666_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_666_inst_ack_1 : boolean;
  signal type_cast_670_inst_req_0 : boolean;
  signal type_cast_670_inst_ack_0 : boolean;
  signal type_cast_670_inst_req_1 : boolean;
  signal type_cast_670_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_684_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_684_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_684_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_684_inst_ack_1 : boolean;
  signal type_cast_688_inst_req_0 : boolean;
  signal type_cast_688_inst_ack_0 : boolean;
  signal type_cast_688_inst_req_1 : boolean;
  signal type_cast_688_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_702_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_702_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_702_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_702_inst_ack_1 : boolean;
  signal type_cast_706_inst_req_0 : boolean;
  signal type_cast_706_inst_ack_0 : boolean;
  signal type_cast_706_inst_req_1 : boolean;
  signal type_cast_706_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_720_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_720_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_720_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_720_inst_ack_1 : boolean;
  signal type_cast_724_inst_req_0 : boolean;
  signal type_cast_724_inst_ack_0 : boolean;
  signal type_cast_724_inst_req_1 : boolean;
  signal type_cast_724_inst_ack_1 : boolean;
  signal ptr_deref_732_store_0_req_0 : boolean;
  signal ptr_deref_732_store_0_ack_0 : boolean;
  signal ptr_deref_732_store_0_req_1 : boolean;
  signal ptr_deref_732_store_0_ack_1 : boolean;
  signal if_stmt_746_branch_req_0 : boolean;
  signal if_stmt_746_branch_ack_1 : boolean;
  signal if_stmt_746_branch_ack_0 : boolean;
  signal type_cast_757_inst_req_0 : boolean;
  signal type_cast_757_inst_ack_0 : boolean;
  signal type_cast_757_inst_req_1 : boolean;
  signal type_cast_757_inst_ack_1 : boolean;
  signal type_cast_338_inst_req_0 : boolean;
  signal type_cast_338_inst_ack_0 : boolean;
  signal type_cast_338_inst_req_1 : boolean;
  signal type_cast_338_inst_ack_1 : boolean;
  signal phi_stmt_335_req_0 : boolean;
  signal type_cast_345_inst_req_0 : boolean;
  signal type_cast_345_inst_ack_0 : boolean;
  signal type_cast_345_inst_req_1 : boolean;
  signal type_cast_345_inst_ack_1 : boolean;
  signal phi_stmt_342_req_0 : boolean;
  signal phi_stmt_335_req_1 : boolean;
  signal type_cast_347_inst_req_0 : boolean;
  signal type_cast_347_inst_ack_0 : boolean;
  signal type_cast_347_inst_req_1 : boolean;
  signal type_cast_347_inst_ack_1 : boolean;
  signal phi_stmt_342_req_1 : boolean;
  signal phi_stmt_335_ack_0 : boolean;
  signal phi_stmt_342_ack_0 : boolean;
  signal type_cast_408_inst_req_0 : boolean;
  signal type_cast_408_inst_ack_0 : boolean;
  signal type_cast_408_inst_req_1 : boolean;
  signal type_cast_408_inst_ack_1 : boolean;
  signal phi_stmt_405_req_0 : boolean;
  signal phi_stmt_405_ack_0 : boolean;
  signal type_cast_415_inst_req_0 : boolean;
  signal type_cast_415_inst_ack_0 : boolean;
  signal type_cast_415_inst_req_1 : boolean;
  signal type_cast_415_inst_ack_1 : boolean;
  signal phi_stmt_412_req_0 : boolean;
  signal type_cast_417_inst_req_0 : boolean;
  signal type_cast_417_inst_ack_0 : boolean;
  signal type_cast_417_inst_req_1 : boolean;
  signal type_cast_417_inst_ack_1 : boolean;
  signal phi_stmt_412_req_1 : boolean;
  signal phi_stmt_412_ack_0 : boolean;
  signal phi_stmt_583_req_0 : boolean;
  signal type_cast_589_inst_req_0 : boolean;
  signal type_cast_589_inst_ack_0 : boolean;
  signal type_cast_589_inst_req_1 : boolean;
  signal type_cast_589_inst_ack_1 : boolean;
  signal phi_stmt_583_req_1 : boolean;
  signal phi_stmt_583_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_684_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_684_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_684_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_684_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_684: Block -- control-path 
    signal testConfigure_CP_684_elements: BooleanArray(291 downto 0);
    -- 
  begin -- 
    testConfigure_CP_684_elements(0) <= testConfigure_CP_684_start;
    testConfigure_CP_684_symbol <= testConfigure_CP_684_elements(256);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	30 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	35 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	38 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	50 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	22 
    -- CP-element group 0: 	24 
    -- CP-element group 0:  members (112) 
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_3_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_3_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_3_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_3_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_2_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_3_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325__entry__
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_1_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_1_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_3_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_3_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_1_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_2_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_0_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_0_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_0_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_3/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_2_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_3/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_2_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_2_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_2_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/branch_block_stmt_275__entry__
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_1_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_2/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_1_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_2/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_0_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_1_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_1_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_1/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_0_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_1_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_0_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_0_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_update_start_
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_0_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_update_start
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_sample_start
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_275/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_addr_resize/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_update_start_
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_update_start_
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_update_start
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_2_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_sample_start
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_2_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_update_start_
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_3_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_1/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_2/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_2/cr
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_3/$entry
      -- CP-element group 0: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_3/cr
      -- 
    cr_1004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_addr_3_req_1); -- 
    rr_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_addr_3_req_0); -- 
    cr_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_297_store_0_req_1); -- 
    rr_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_addr_1_req_0); -- 
    rr_859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => RPIPE_zeropad_input_pipe_288_inst_req_0); -- 
    cr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_305_inst_req_1); -- 
    rr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_addr_3_req_0); -- 
    cr_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_addr_1_req_1); -- 
    cr_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_addr_2_req_1); -- 
    cr_974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_addr_0_req_1); -- 
    cr_850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_store_3_req_1); -- 
    rr_778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_addr_2_req_0); -- 
    cr_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_addr_2_req_1); -- 
    cr_773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_addr_1_req_1); -- 
    cr_845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_store_2_req_1); -- 
    rr_969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_addr_0_req_0); -- 
    rr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_addr_1_req_0); -- 
    cr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_store_1_req_1); -- 
    cr_835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_store_0_req_1); -- 
    cr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_addr_0_req_1); -- 
    rr_758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_addr_0_req_0); -- 
    rr_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_addr_2_req_0); -- 
    cr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_283_addr_3_req_1); -- 
    cr_1046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_store_0_req_1); -- 
    cr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_store_1_req_1); -- 
    cr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_store_2_req_1); -- 
    cr_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_314_store_3_req_1); -- 
    -- CP-element group 1:  join  fork  transition  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: 	3 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	12 
    -- CP-element group 1: 	13 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	15 
    -- CP-element group 1:  members (15) 
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_0/rr
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_0/$entry
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/$entry
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/ptr_deref_283_Split/split_ack
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/ptr_deref_283_Split/split_req
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/ptr_deref_283_Split/$exit
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/ptr_deref_283_Split/$entry
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_3/rr
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_3/$entry
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_2/rr
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_2/$entry
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_1/rr
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_1/$entry
      -- CP-element group 1: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_sample_start_
      -- 
    rr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(1), ack => ptr_deref_283_store_0_req_0); -- 
    rr_814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(1), ack => ptr_deref_283_store_1_req_0); -- 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(1), ack => ptr_deref_283_store_2_req_0); -- 
    rr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(1), ack => ptr_deref_283_store_3_req_0); -- 
    testConfigure_cp_element_group_1: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_1"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(0) & testConfigure_CP_684_elements(3);
      gj_testConfigure_cp_element_group_1 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(1), clk => clk, reset => reset); --
    end block;
    -- CP-element group 2:  join  transition  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	56 
    -- CP-element group 2:  members (1) 
      -- CP-element group 2: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_sample_complete
      -- 
    testConfigure_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(4) & testConfigure_CP_684_elements(6) & testConfigure_CP_684_elements(8) & testConfigure_CP_684_elements(10);
      gj_testConfigure_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	7 
    -- CP-element group 3: 	9 
    -- CP-element group 3: 	11 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	1 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_update_complete
      -- CP-element group 3: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_address_calculated
      -- 
    testConfigure_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(5) & testConfigure_CP_684_elements(7) & testConfigure_CP_684_elements(9) & testConfigure_CP_684_elements(11);
      gj_testConfigure_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	2 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_0_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_0_Sample/$exit
      -- 
    ra_759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_addr_0_ack_0, ack => testConfigure_CP_684_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	3 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_0_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_0_Update/$exit
      -- 
    ca_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_addr_0_ack_1, ack => testConfigure_CP_684_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	2 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_1_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_1_Sample/$exit
      -- 
    ra_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_addr_1_ack_0, ack => testConfigure_CP_684_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	3 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_1_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_1_Update/$exit
      -- 
    ca_774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_addr_1_ack_1, ack => testConfigure_CP_684_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_2_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_2_Sample/$exit
      -- 
    ra_779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_addr_2_ack_0, ack => testConfigure_CP_684_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	3 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_2_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_2_Update/$exit
      -- 
    ca_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_addr_2_ack_1, ack => testConfigure_CP_684_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	2 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_3_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_3_Sample/$exit
      -- 
    ra_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_addr_3_ack_0, ack => testConfigure_CP_684_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	3 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_3_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_word_addrgen_3_Update/ca
      -- 
    ca_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_addr_3_ack_1, ack => testConfigure_CP_684_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	1 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_0/ra
      -- 
    ra_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_store_0_ack_0, ack => testConfigure_CP_684_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	1 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_1/ra
      -- CP-element group 13: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_1/$exit
      -- 
    ra_815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_store_1_ack_0, ack => testConfigure_CP_684_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_2/ra
      -- CP-element group 14: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_2/$exit
      -- 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_store_2_ack_0, ack => testConfigure_CP_684_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	1 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_3/$exit
      -- CP-element group 15: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/word_3/ra
      -- 
    ra_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_store_3_ack_0, ack => testConfigure_CP_684_elements(15)); -- 
    -- CP-element group 16:  join  transition  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: 	13 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	54 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_sample_completed_
      -- 
    testConfigure_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(12) & testConfigure_CP_684_elements(13) & testConfigure_CP_684_elements(14) & testConfigure_CP_684_elements(15);
      gj_testConfigure_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	21 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_0/$exit
      -- 
    ca_836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_store_0_ack_1, ack => testConfigure_CP_684_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_1/ca
      -- CP-element group 18: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_1/$exit
      -- 
    ca_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_store_1_ack_1, ack => testConfigure_CP_684_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_2/ca
      -- CP-element group 19: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_2/$exit
      -- 
    ca_846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_store_2_ack_1, ack => testConfigure_CP_684_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_3/ca
      -- CP-element group 20: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/word_3/$exit
      -- 
    ca_851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_283_store_3_ack_1, ack => testConfigure_CP_684_elements(20)); -- 
    -- CP-element group 21:  join  transition  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	19 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	56 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_update_completed_
      -- 
    testConfigure_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(17) & testConfigure_CP_684_elements(18) & testConfigure_CP_684_elements(19) & testConfigure_CP_684_elements(20);
      gj_testConfigure_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	0 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_update_start_
      -- CP-element group 22: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_sample_completed_
      -- 
    ra_860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_288_inst_ack_0, ack => testConfigure_CP_684_elements(22)); -- 
    cr_864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(22), ack => RPIPE_zeropad_input_pipe_288_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_288_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_sample_start_
      -- 
    ca_865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_288_inst_ack_1, ack => testConfigure_CP_684_elements(23)); -- 
    rr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(23), ack => RPIPE_zeropad_input_pipe_301_inst_req_0); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: 	54 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/ptr_deref_297_Split/$exit
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/ptr_deref_297_Split/$entry
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/word_access_start/word_0/rr
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/word_access_start/word_0/$entry
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/word_access_start/$entry
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/ptr_deref_297_Split/split_ack
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/ptr_deref_297_Split/split_req
      -- CP-element group 24: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_sample_start_
      -- 
    rr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(24), ack => ptr_deref_297_store_0_req_0); -- 
    testConfigure_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(0) & testConfigure_CP_684_elements(54) & testConfigure_CP_684_elements(23);
      gj_testConfigure_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	55 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_sample_completed_
      -- 
    ra_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_297_store_0_ack_0, ack => testConfigure_CP_684_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	56 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_update_completed_
      -- 
    ca_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_297_store_0_ack_1, ack => testConfigure_CP_684_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_update_start_
      -- CP-element group 27: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_sample_completed_
      -- 
    ra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_301_inst_ack_0, ack => testConfigure_CP_684_elements(27)); -- 
    cr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(27), ack => RPIPE_zeropad_input_pipe_301_inst_req_1); -- 
    -- CP-element group 28:  fork  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	52 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_301_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_Sample/rr
      -- 
    ca_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_301_inst_ack_1, ack => testConfigure_CP_684_elements(28)); -- 
    rr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(28), ack => type_cast_305_inst_req_0); -- 
    rr_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(28), ack => RPIPE_zeropad_input_pipe_324_inst_req_0); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_Sample/$exit
      -- 
    ra_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_0, ack => testConfigure_CP_684_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	0 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/type_cast_305_update_completed_
      -- 
    ca_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_1, ack => testConfigure_CP_684_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	55 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	42 
    -- CP-element group 31: 	43 
    -- CP-element group 31: 	44 
    -- CP-element group 31: 	45 
    -- CP-element group 31:  members (15) 
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/ptr_deref_314_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/ptr_deref_314_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/ptr_deref_314_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/ptr_deref_314_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_0/rr
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_1/$entry
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_1/rr
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_2/$entry
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_2/rr
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_3/$entry
      -- CP-element group 31: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_3/rr
      -- 
    rr_1020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(31), ack => ptr_deref_314_store_0_req_0); -- 
    rr_1025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(31), ack => ptr_deref_314_store_1_req_0); -- 
    rr_1030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(31), ack => ptr_deref_314_store_2_req_0); -- 
    rr_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(31), ack => ptr_deref_314_store_3_req_0); -- 
    testConfigure_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(0) & testConfigure_CP_684_elements(30) & testConfigure_CP_684_elements(33) & testConfigure_CP_684_elements(55);
      gj_testConfigure_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: 	36 
    -- CP-element group 32: 	38 
    -- CP-element group 32: 	40 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	56 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_sample_complete
      -- 
    testConfigure_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(34) & testConfigure_CP_684_elements(36) & testConfigure_CP_684_elements(38) & testConfigure_CP_684_elements(40);
      gj_testConfigure_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: 	37 
    -- CP-element group 33: 	39 
    -- CP-element group 33: 	41 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_update_complete
      -- 
    testConfigure_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(35) & testConfigure_CP_684_elements(37) & testConfigure_CP_684_elements(39) & testConfigure_CP_684_elements(41);
      gj_testConfigure_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_0_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_0_Sample/$exit
      -- 
    ra_970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_addr_0_ack_0, ack => testConfigure_CP_684_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	0 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_0_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_0_Update/$exit
      -- 
    ca_975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_addr_0_ack_1, ack => testConfigure_CP_684_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	32 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_1_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_1_Sample/ra
      -- 
    ra_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_addr_1_ack_0, ack => testConfigure_CP_684_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	33 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_1_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_1_Update/ca
      -- 
    ca_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_addr_1_ack_1, ack => testConfigure_CP_684_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	0 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_2_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_2_Sample/$exit
      -- 
    ra_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_addr_2_ack_0, ack => testConfigure_CP_684_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	33 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_2_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_2_Update/$exit
      -- 
    ca_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_addr_2_ack_1, ack => testConfigure_CP_684_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	32 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_3_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_3_Sample/ra
      -- 
    ra_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_addr_3_ack_0, ack => testConfigure_CP_684_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	33 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_3_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_word_addrgen_3_Update/ca
      -- 
    ca_1005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_addr_3_ack_1, ack => testConfigure_CP_684_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	31 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	46 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_0/ra
      -- 
    ra_1021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_store_0_ack_0, ack => testConfigure_CP_684_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	31 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_1/ra
      -- 
    ra_1026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_store_1_ack_0, ack => testConfigure_CP_684_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	31 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_2/$exit
      -- CP-element group 44: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_2/ra
      -- 
    ra_1031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_store_2_ack_0, ack => testConfigure_CP_684_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	31 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_3/$exit
      -- CP-element group 45: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/word_3/ra
      -- 
    ra_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_store_3_ack_0, ack => testConfigure_CP_684_elements(45)); -- 
    -- CP-element group 46:  join  transition  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	42 
    -- CP-element group 46: 	43 
    -- CP-element group 46: 	44 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/word_access_start/$exit
      -- CP-element group 46: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_sample_completed_
      -- 
    testConfigure_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(42) & testConfigure_CP_684_elements(43) & testConfigure_CP_684_elements(44) & testConfigure_CP_684_elements(45);
      gj_testConfigure_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	51 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_0/ca
      -- 
    ca_1047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_store_0_ack_1, ack => testConfigure_CP_684_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	51 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_1/ca
      -- 
    ca_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_store_1_ack_1, ack => testConfigure_CP_684_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_2/$exit
      -- CP-element group 49: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_2/ca
      -- 
    ca_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_store_2_ack_1, ack => testConfigure_CP_684_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	0 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_3/$exit
      -- CP-element group 50: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/word_3/ca
      -- 
    ca_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_314_store_3_ack_1, ack => testConfigure_CP_684_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	47 
    -- CP-element group 51: 	48 
    -- CP-element group 51: 	49 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	56 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_314_Update/word_access_complete/$exit
      -- 
    testConfigure_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(47) & testConfigure_CP_684_elements(48) & testConfigure_CP_684_elements(49) & testConfigure_CP_684_elements(50);
      gj_testConfigure_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	28 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_update_start_
      -- CP-element group 52: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_Update/cr
      -- 
    ra_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_324_inst_ack_0, ack => testConfigure_CP_684_elements(52)); -- 
    cr_1075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(52), ack => RPIPE_zeropad_input_pipe_324_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/RPIPE_zeropad_input_pipe_324_Update/ca
      -- 
    ca_1076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_324_inst_ack_1, ack => testConfigure_CP_684_elements(53)); -- 
    -- CP-element group 54:  transition  delay-element  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	16 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	24 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_283_ptr_deref_297_delay
      -- 
    -- Element group testConfigure_CP_684_elements(54) is a control-delay.
    cp_element_54_delay: control_delay_element  generic map(name => " 54_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(16), ack => testConfigure_CP_684_elements(54), clk => clk, reset =>reset);
    -- CP-element group 55:  transition  delay-element  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	25 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	31 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/ptr_deref_297_ptr_deref_314_delay
      -- 
    -- Element group testConfigure_CP_684_elements(55) is a control-delay.
    cp_element_55_delay: control_delay_element  generic map(name => " 55_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(25), ack => testConfigure_CP_684_elements(55), clk => clk, reset =>reset);
    -- CP-element group 56:  branch  join  transition  place  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	26 
    -- CP-element group 56: 	32 
    -- CP-element group 56: 	51 
    -- CP-element group 56: 	53 
    -- CP-element group 56: 	2 
    -- CP-element group 56: 	21 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (10) 
      -- CP-element group 56: 	 branch_block_stmt_275/if_stmt_326__entry__
      -- CP-element group 56: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325__exit__
      -- CP-element group 56: 	 branch_block_stmt_275/assign_stmt_281_to_assign_stmt_325/$exit
      -- CP-element group 56: 	 branch_block_stmt_275/if_stmt_326_dead_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_275/if_stmt_326_eval_test/$entry
      -- CP-element group 56: 	 branch_block_stmt_275/if_stmt_326_eval_test/$exit
      -- CP-element group 56: 	 branch_block_stmt_275/if_stmt_326_eval_test/branch_req
      -- CP-element group 56: 	 branch_block_stmt_275/R_cmp86_327_place
      -- CP-element group 56: 	 branch_block_stmt_275/if_stmt_326_if_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_275/if_stmt_326_else_link/$entry
      -- 
    branch_req_1086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(56), ack => if_stmt_326_branch_req_0); -- 
    testConfigure_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(26) & testConfigure_CP_684_elements(32) & testConfigure_CP_684_elements(51) & testConfigure_CP_684_elements(53) & testConfigure_CP_684_elements(2) & testConfigure_CP_684_elements(21);
      gj_testConfigure_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	277 
    -- CP-element group 57: 	278 
    -- CP-element group 57:  members (12) 
      -- CP-element group 57: 	 branch_block_stmt_275/if_stmt_326_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_275/if_stmt_326_if_link/if_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/$entry
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/$entry
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/$entry
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/$entry
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/Update/cr
      -- 
    if_choice_transition_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_326_branch_ack_1, ack => testConfigure_CP_684_elements(57)); -- 
    rr_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(57), ack => type_cast_415_inst_req_0); -- 
    cr_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(57), ack => type_cast_415_inst_req_1); -- 
    -- CP-element group 58:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	264 
    -- CP-element group 58: 	265 
    -- CP-element group 58: 	266 
    -- CP-element group 58:  members (22) 
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 58: 	 branch_block_stmt_275/merge_stmt_332__exit__
      -- CP-element group 58: 	 branch_block_stmt_275/if_stmt_326_else_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_275/if_stmt_326_else_link/else_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_275/entry_forx_xbodyx_xpreheader
      -- CP-element group 58: 	 branch_block_stmt_275/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_275/merge_stmt_332_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_275/merge_stmt_332_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/merge_stmt_332_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_275/merge_stmt_332_PhiAck/dummy
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_335/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_326_branch_ack_0, ack => testConfigure_CP_684_elements(58)); -- 
    rr_2581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(58), ack => type_cast_347_inst_req_0); -- 
    cr_2586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(58), ack => type_cast_347_inst_req_1); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	272 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_Sample/ra
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_0, ack => testConfigure_CP_684_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	272 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	114 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_Update/ca
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_1, ack => testConfigure_CP_684_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	272 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	114 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_sample_complete
      -- CP-element group 61: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_Sample/ra
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_363_index_1_scale_ack_0, ack => testConfigure_CP_684_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	272 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scaled_1
      -- CP-element group 62: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_update_complete
      -- CP-element group 62: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_Sample/req
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_363_index_1_scale_ack_1, ack => testConfigure_CP_684_elements(62)); -- 
    req_1148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(62), ack => array_obj_ref_363_index_offset_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	114 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_sample_complete
      -- CP-element group 63: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_Sample/ack
      -- 
    ack_1149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_363_index_offset_ack_0, ack => testConfigure_CP_684_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	272 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (11) 
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_root_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_offset_calculated
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_base_plus_offset/$entry
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_base_plus_offset/$exit
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_base_plus_offset/sum_rename_req
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_base_plus_offset/sum_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_request/$entry
      -- CP-element group 64: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_request/req
      -- 
    ack_1154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_363_index_offset_ack_1, ack => testConfigure_CP_684_elements(64)); -- 
    req_1163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(64), ack => addr_of_364_final_reg_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_request/$exit
      -- CP-element group 65: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_request/ack
      -- 
    ack_1164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_364_final_reg_ack_0, ack => testConfigure_CP_684_elements(65)); -- 
    -- CP-element group 66:  fork  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	272 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	69 
    -- CP-element group 66: 	72 
    -- CP-element group 66: 	74 
    -- CP-element group 66: 	76 
    -- CP-element group 66: 	78 
    -- CP-element group 66:  members (23) 
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_complete/ack
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_address_calculated
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_root_address_calculated
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_address_resized
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_addr_resize/$entry
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_addr_resize/$exit
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_addr_resize/base_resize_req
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_addr_resize/base_resize_ack
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_plus_offset/$entry
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_plus_offset/$exit
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_plus_offset/sum_rename_req
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_base_plus_offset/sum_rename_ack
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_sample_start
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_0_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_0_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_1_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_1_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_2_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_2_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_3_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_3_Sample/rr
      -- 
    ack_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_364_final_reg_ack_1, ack => testConfigure_CP_684_elements(66)); -- 
    rr_1209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(66), ack => ptr_deref_371_addr_0_req_0); -- 
    rr_1219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(66), ack => ptr_deref_371_addr_1_req_0); -- 
    rr_1229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(66), ack => ptr_deref_371_addr_2_req_0); -- 
    rr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(66), ack => ptr_deref_371_addr_3_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	272 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_Sample/ra
      -- 
    ra_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_368_inst_ack_0, ack => testConfigure_CP_684_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	272 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_Update/ca
      -- 
    ca_1183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_368_inst_ack_1, ack => testConfigure_CP_684_elements(68)); -- 
    -- CP-element group 69:  join  fork  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	66 
    -- CP-element group 69: 	68 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	80 
    -- CP-element group 69: 	81 
    -- CP-element group 69: 	82 
    -- CP-element group 69: 	83 
    -- CP-element group 69:  members (15) 
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/ptr_deref_371_Split/$entry
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/ptr_deref_371_Split/$exit
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/ptr_deref_371_Split/split_req
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/ptr_deref_371_Split/split_ack
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/$entry
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_0/$entry
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_0/rr
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_1/$entry
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_1/rr
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_2/$entry
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_2/rr
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_3/$entry
      -- CP-element group 69: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_3/rr
      -- 
    rr_1260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(69), ack => ptr_deref_371_store_0_req_0); -- 
    rr_1265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(69), ack => ptr_deref_371_store_1_req_0); -- 
    rr_1270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(69), ack => ptr_deref_371_store_2_req_0); -- 
    rr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(69), ack => ptr_deref_371_store_3_req_0); -- 
    testConfigure_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(66) & testConfigure_CP_684_elements(68) & testConfigure_CP_684_elements(71);
      gj_testConfigure_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70: 	76 
    -- CP-element group 70: 	78 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	114 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_sample_complete
      -- 
    testConfigure_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(72) & testConfigure_CP_684_elements(74) & testConfigure_CP_684_elements(76) & testConfigure_CP_684_elements(78);
      gj_testConfigure_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	75 
    -- CP-element group 71: 	77 
    -- CP-element group 71: 	79 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_address_calculated
      -- CP-element group 71: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_update_complete
      -- 
    testConfigure_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(73) & testConfigure_CP_684_elements(75) & testConfigure_CP_684_elements(77) & testConfigure_CP_684_elements(79);
      gj_testConfigure_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	66 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_0_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_0_Sample/ra
      -- 
    ra_1210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_addr_0_ack_0, ack => testConfigure_CP_684_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	272 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_0_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_0_Update/ca
      -- 
    ca_1215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_addr_0_ack_1, ack => testConfigure_CP_684_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	66 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	70 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_1_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_1_Sample/ra
      -- 
    ra_1220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_addr_1_ack_0, ack => testConfigure_CP_684_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	272 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	71 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_1_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_1_Update/ca
      -- 
    ca_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_addr_1_ack_1, ack => testConfigure_CP_684_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	66 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	70 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_2_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_2_Sample/ra
      -- 
    ra_1230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_addr_2_ack_0, ack => testConfigure_CP_684_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	272 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	71 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_2_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_2_Update/ca
      -- 
    ca_1235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_addr_2_ack_1, ack => testConfigure_CP_684_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	66 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	70 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_3_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_3_Sample/ra
      -- 
    ra_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_addr_3_ack_0, ack => testConfigure_CP_684_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	272 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	71 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_3_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_3_Update/ca
      -- 
    ca_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_addr_3_ack_1, ack => testConfigure_CP_684_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	69 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	84 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_0/ra
      -- 
    ra_1261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_store_0_ack_0, ack => testConfigure_CP_684_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	69 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	84 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_1/$exit
      -- CP-element group 81: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_1/ra
      -- 
    ra_1266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_store_1_ack_0, ack => testConfigure_CP_684_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	69 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_2/$exit
      -- CP-element group 82: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_2/ra
      -- 
    ra_1271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_store_2_ack_0, ack => testConfigure_CP_684_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	69 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_3/$exit
      -- CP-element group 83: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/word_3/ra
      -- 
    ra_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_store_3_ack_0, ack => testConfigure_CP_684_elements(83)); -- 
    -- CP-element group 84:  join  transition  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: 	81 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	113 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Sample/word_access_start/$exit
      -- 
    testConfigure_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(80) & testConfigure_CP_684_elements(81) & testConfigure_CP_684_elements(82) & testConfigure_CP_684_elements(83);
      gj_testConfigure_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	272 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	89 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_0/ca
      -- 
    ca_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_store_0_ack_1, ack => testConfigure_CP_684_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	272 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	89 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_1/$exit
      -- CP-element group 86: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_1/ca
      -- 
    ca_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_store_1_ack_1, ack => testConfigure_CP_684_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	272 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_2/$exit
      -- CP-element group 87: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_2/ca
      -- 
    ca_1297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_store_2_ack_1, ack => testConfigure_CP_684_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	272 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_3/$exit
      -- CP-element group 88: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_3/ca
      -- 
    ca_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_371_store_3_ack_1, ack => testConfigure_CP_684_elements(88)); -- 
    -- CP-element group 89:  join  transition  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	85 
    -- CP-element group 89: 	86 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	114 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/$exit
      -- 
    testConfigure_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(85) & testConfigure_CP_684_elements(86) & testConfigure_CP_684_elements(87) & testConfigure_CP_684_elements(88);
      gj_testConfigure_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  fork  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: 	113 
    -- CP-element group 90: 	272 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	101 
    -- CP-element group 90: 	102 
    -- CP-element group 90: 	103 
    -- CP-element group 90: 	104 
    -- CP-element group 90:  members (11) 
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/$entry
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_0/$entry
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_0/rr
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_1/$entry
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_1/rr
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_2/$entry
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_2/rr
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_3/$entry
      -- CP-element group 90: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_3/rr
      -- 
    rr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(90), ack => ptr_deref_388_load_0_req_0); -- 
    rr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(90), ack => ptr_deref_388_load_1_req_0); -- 
    rr_1384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(90), ack => ptr_deref_388_load_2_req_0); -- 
    rr_1389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(90), ack => ptr_deref_388_load_3_req_0); -- 
    testConfigure_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(92) & testConfigure_CP_684_elements(113) & testConfigure_CP_684_elements(272);
      gj_testConfigure_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  transition  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: 	95 
    -- CP-element group 91: 	97 
    -- CP-element group 91: 	99 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	114 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_sample_complete
      -- 
    testConfigure_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(93) & testConfigure_CP_684_elements(95) & testConfigure_CP_684_elements(97) & testConfigure_CP_684_elements(99);
      gj_testConfigure_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: 	96 
    -- CP-element group 92: 	98 
    -- CP-element group 92: 	100 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_address_calculated
      -- CP-element group 92: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_update_complete
      -- 
    testConfigure_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(94) & testConfigure_CP_684_elements(96) & testConfigure_CP_684_elements(98) & testConfigure_CP_684_elements(100);
      gj_testConfigure_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	272 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_0_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_0_Sample/ra
      -- 
    ra_1329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_addr_0_ack_0, ack => testConfigure_CP_684_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	272 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_0_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_0_Update/ca
      -- 
    ca_1334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_addr_0_ack_1, ack => testConfigure_CP_684_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	272 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	91 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_1_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_1_Sample/ra
      -- 
    ra_1339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_addr_1_ack_0, ack => testConfigure_CP_684_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	272 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	92 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_1_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_1_Update/ca
      -- 
    ca_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_addr_1_ack_1, ack => testConfigure_CP_684_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	272 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	91 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_2_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_2_Sample/ra
      -- 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_addr_2_ack_0, ack => testConfigure_CP_684_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	272 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	92 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_2_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_2_Update/ca
      -- 
    ca_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_addr_2_ack_1, ack => testConfigure_CP_684_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	272 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	91 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_3_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_3_Sample/ra
      -- 
    ra_1359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_addr_3_ack_0, ack => testConfigure_CP_684_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	272 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	92 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_3_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_3_Update/ca
      -- 
    ca_1364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_addr_3_ack_1, ack => testConfigure_CP_684_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	90 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	105 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_0/ra
      -- 
    ra_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_load_0_ack_0, ack => testConfigure_CP_684_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	90 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	105 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_1/$exit
      -- CP-element group 102: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_1/ra
      -- 
    ra_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_load_1_ack_0, ack => testConfigure_CP_684_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	90 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_2/$exit
      -- CP-element group 103: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_2/ra
      -- 
    ra_1385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_load_2_ack_0, ack => testConfigure_CP_684_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	90 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_3/$exit
      -- CP-element group 104: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/word_3/ra
      -- 
    ra_1390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_load_3_ack_0, ack => testConfigure_CP_684_elements(104)); -- 
    -- CP-element group 105:  join  transition  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	101 
    -- CP-element group 105: 	102 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Sample/word_access_start/$exit
      -- 
    testConfigure_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(101) & testConfigure_CP_684_elements(102) & testConfigure_CP_684_elements(103) & testConfigure_CP_684_elements(104);
      gj_testConfigure_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	272 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_0/$exit
      -- CP-element group 106: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_0/ca
      -- 
    ca_1401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_load_0_ack_1, ack => testConfigure_CP_684_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	272 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_1/$exit
      -- CP-element group 107: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_1/ca
      -- 
    ca_1406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_load_1_ack_1, ack => testConfigure_CP_684_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	272 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_2/$exit
      -- CP-element group 108: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_2/ca
      -- 
    ca_1411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_load_2_ack_1, ack => testConfigure_CP_684_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	272 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_3/$exit
      -- CP-element group 109: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_3/ca
      -- 
    ca_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_388_load_3_ack_1, ack => testConfigure_CP_684_elements(109)); -- 
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	106 
    -- CP-element group 110: 	107 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	114 
    -- CP-element group 110:  members (7) 
      -- CP-element group 110: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/ptr_deref_388_Merge/$entry
      -- CP-element group 110: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/ptr_deref_388_Merge/$exit
      -- CP-element group 110: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/ptr_deref_388_Merge/merge_req
      -- CP-element group 110: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/ptr_deref_388_Merge/merge_ack
      -- 
    testConfigure_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(106) & testConfigure_CP_684_elements(107) & testConfigure_CP_684_elements(108) & testConfigure_CP_684_elements(109);
      gj_testConfigure_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	272 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_update_start_
      -- CP-element group 111: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_Update/cr
      -- 
    ra_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_396_inst_ack_0, ack => testConfigure_CP_684_elements(111)); -- 
    cr_1434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(111), ack => RPIPE_zeropad_input_pipe_396_inst_req_1); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_Update/ca
      -- 
    ca_1435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_396_inst_ack_1, ack => testConfigure_CP_684_elements(112)); -- 
    -- CP-element group 113:  transition  delay-element  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	84 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	90 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_ptr_deref_388_delay
      -- 
    -- Element group testConfigure_CP_684_elements(113) is a control-delay.
    cp_element_113_delay: control_delay_element  generic map(name => " 113_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(84), ack => testConfigure_CP_684_elements(113), clk => clk, reset =>reset);
    -- CP-element group 114:  branch  join  transition  place  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	70 
    -- CP-element group 114: 	89 
    -- CP-element group 114: 	91 
    -- CP-element group 114: 	60 
    -- CP-element group 114: 	61 
    -- CP-element group 114: 	63 
    -- CP-element group 114: 	110 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (10) 
      -- CP-element group 114: 	 branch_block_stmt_275/if_stmt_398__entry__
      -- CP-element group 114: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397__exit__
      -- CP-element group 114: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/$exit
      -- CP-element group 114: 	 branch_block_stmt_275/if_stmt_398_dead_link/$entry
      -- CP-element group 114: 	 branch_block_stmt_275/if_stmt_398_eval_test/$entry
      -- CP-element group 114: 	 branch_block_stmt_275/if_stmt_398_eval_test/$exit
      -- CP-element group 114: 	 branch_block_stmt_275/if_stmt_398_eval_test/branch_req
      -- CP-element group 114: 	 branch_block_stmt_275/R_cmp_399_place
      -- CP-element group 114: 	 branch_block_stmt_275/if_stmt_398_if_link/$entry
      -- CP-element group 114: 	 branch_block_stmt_275/if_stmt_398_else_link/$entry
      -- 
    branch_req_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(114), ack => if_stmt_398_branch_req_0); -- 
    testConfigure_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(70) & testConfigure_CP_684_elements(89) & testConfigure_CP_684_elements(91) & testConfigure_CP_684_elements(60) & testConfigure_CP_684_elements(61) & testConfigure_CP_684_elements(63) & testConfigure_CP_684_elements(110) & testConfigure_CP_684_elements(112);
      gj_testConfigure_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  place  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	257 
    -- CP-element group 115: 	258 
    -- CP-element group 115: 	260 
    -- CP-element group 115: 	261 
    -- CP-element group 115:  members (20) 
      -- CP-element group 115: 	 branch_block_stmt_275/if_stmt_398_if_link/$exit
      -- CP-element group 115: 	 branch_block_stmt_275/if_stmt_398_if_link/if_choice_transition
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/Update/cr
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/Update/cr
      -- 
    if_choice_transition_1449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_398_branch_ack_1, ack => testConfigure_CP_684_elements(115)); -- 
    rr_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(115), ack => type_cast_338_inst_req_0); -- 
    cr_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(115), ack => type_cast_338_inst_req_1); -- 
    rr_2547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(115), ack => type_cast_345_inst_req_0); -- 
    cr_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(115), ack => type_cast_345_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  place  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	273 
    -- CP-element group 116: 	274 
    -- CP-element group 116:  members (12) 
      -- CP-element group 116: 	 branch_block_stmt_275/if_stmt_398_else_link/$exit
      -- CP-element group 116: 	 branch_block_stmt_275/if_stmt_398_else_link/else_choice_transition
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/$entry
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/$entry
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/$entry
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/$entry
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_398_branch_ack_0, ack => testConfigure_CP_684_elements(116)); -- 
    rr_2617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(116), ack => type_cast_408_inst_req_0); -- 
    cr_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(116), ack => type_cast_408_inst_req_1); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	284 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/word_access_start/word_0/ra
      -- 
    ra_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_419_store_0_ack_0, ack => testConfigure_CP_684_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	284 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	208 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Update/word_access_complete/word_0/ca
      -- 
    ca_1491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_419_store_0_ack_1, ack => testConfigure_CP_684_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	284 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_update_start_
      -- CP-element group 119: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_Update/cr
      -- 
    ra_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_423_inst_ack_0, ack => testConfigure_CP_684_elements(119)); -- 
    cr_1504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(119), ack => RPIPE_zeropad_input_pipe_423_inst_req_1); -- 
    -- CP-element group 120:  fork  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: 	126 
    -- CP-element group 120:  members (9) 
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_Sample/rr
      -- 
    ca_1505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_423_inst_ack_1, ack => testConfigure_CP_684_elements(120)); -- 
    rr_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(120), ack => type_cast_427_inst_req_0); -- 
    rr_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(120), ack => RPIPE_zeropad_input_pipe_442_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_Sample/ra
      -- 
    ra_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_427_inst_ack_0, ack => testConfigure_CP_684_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	284 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_Update/ca
      -- 
    ca_1519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_427_inst_ack_1, ack => testConfigure_CP_684_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: 	284 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/ptr_deref_438_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/ptr_deref_438_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/ptr_deref_438_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/ptr_deref_438_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/word_access_start/word_0/rr
      -- 
    rr_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(123), ack => ptr_deref_438_store_0_req_0); -- 
    testConfigure_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(122) & testConfigure_CP_684_elements(284);
      gj_testConfigure_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	206 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Sample/word_access_start/word_0/ra
      -- 
    ra_1558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_438_store_0_ack_0, ack => testConfigure_CP_684_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	284 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	208 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Update/word_access_complete/word_0/ca
      -- 
    ca_1569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_438_store_0_ack_1, ack => testConfigure_CP_684_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	120 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_update_start_
      -- CP-element group 126: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_Sample/ra
      -- CP-element group 126: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_Update/cr
      -- 
    ra_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_442_inst_ack_0, ack => testConfigure_CP_684_elements(126)); -- 
    cr_1582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(126), ack => RPIPE_zeropad_input_pipe_442_inst_req_1); -- 
    -- CP-element group 127:  fork  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: 	133 
    -- CP-element group 127:  members (9) 
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_442_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_Sample/rr
      -- 
    ca_1583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_442_inst_ack_1, ack => testConfigure_CP_684_elements(127)); -- 
    rr_1591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(127), ack => type_cast_446_inst_req_0); -- 
    rr_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(127), ack => RPIPE_zeropad_input_pipe_461_inst_req_0); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_Sample/ra
      -- 
    ra_1592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_446_inst_ack_0, ack => testConfigure_CP_684_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	284 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_Update/ca
      -- 
    ca_1597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_446_inst_ack_1, ack => testConfigure_CP_684_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: 	206 
    -- CP-element group 130: 	284 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/word_access_start/word_0/$entry
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/word_access_start/word_0/rr
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/ptr_deref_457_Split/$entry
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/ptr_deref_457_Split/$exit
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/ptr_deref_457_Split/split_req
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/ptr_deref_457_Split/split_ack
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/word_access_start/$entry
      -- CP-element group 130: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_sample_start_
      -- 
    rr_1635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(130), ack => ptr_deref_457_store_0_req_0); -- 
    testConfigure_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(129) & testConfigure_CP_684_elements(206) & testConfigure_CP_684_elements(284);
      gj_testConfigure_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	207 
    -- CP-element group 131:  members (5) 
      -- CP-element group 131: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/word_access_start/word_0/ra
      -- CP-element group 131: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/word_access_start/word_0/$exit
      -- CP-element group 131: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Sample/word_access_start/$exit
      -- CP-element group 131: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_sample_completed_
      -- 
    ra_1636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_457_store_0_ack_0, ack => testConfigure_CP_684_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	284 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	208 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Update/word_access_complete/$exit
      -- CP-element group 132: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Update/word_access_complete/word_0/$exit
      -- CP-element group 132: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Update/word_access_complete/word_0/ca
      -- CP-element group 132: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_update_completed_
      -- 
    ca_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_457_store_0_ack_1, ack => testConfigure_CP_684_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	127 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_update_start_
      -- CP-element group 133: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_Sample/$exit
      -- 
    ra_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_461_inst_ack_0, ack => testConfigure_CP_684_elements(133)); -- 
    cr_1660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(133), ack => RPIPE_zeropad_input_pipe_461_inst_req_1); -- 
    -- CP-element group 134:  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_461_Update/$exit
      -- 
    ca_1661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_461_inst_ack_1, ack => testConfigure_CP_684_elements(134)); -- 
    rr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(134), ack => type_cast_465_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_sample_completed_
      -- 
    ra_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_465_inst_ack_0, ack => testConfigure_CP_684_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	284 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_update_completed_
      -- 
    ca_1675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_465_inst_ack_1, ack => testConfigure_CP_684_elements(136)); -- 
    -- CP-element group 137:  join  transition  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: 	207 
    -- CP-element group 137: 	284 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (9) 
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/word_access_start/word_0/$entry
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/ptr_deref_476_Split/$entry
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/ptr_deref_476_Split/$exit
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/ptr_deref_476_Split/split_req
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/ptr_deref_476_Split/split_ack
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/word_access_start/$entry
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/word_access_start/word_0/rr
      -- CP-element group 137: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_sample_start_
      -- 
    rr_1713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(137), ack => ptr_deref_476_store_0_req_0); -- 
    testConfigure_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(136) & testConfigure_CP_684_elements(207) & testConfigure_CP_684_elements(284);
      gj_testConfigure_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (5) 
      -- CP-element group 138: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/word_access_start/$exit
      -- CP-element group 138: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/word_access_start/word_0/$exit
      -- CP-element group 138: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Sample/word_access_start/word_0/ra
      -- CP-element group 138: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_sample_completed_
      -- 
    ra_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_476_store_0_ack_0, ack => testConfigure_CP_684_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	284 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	208 
    -- CP-element group 139:  members (5) 
      -- CP-element group 139: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Update/word_access_complete/$exit
      -- CP-element group 139: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Update/word_access_complete/word_0/$exit
      -- CP-element group 139: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Update/word_access_complete/word_0/ca
      -- CP-element group 139: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_update_completed_
      -- 
    ca_1725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_476_store_0_ack_1, ack => testConfigure_CP_684_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: 	284 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	151 
    -- CP-element group 140: 	152 
    -- CP-element group 140: 	153 
    -- CP-element group 140: 	154 
    -- CP-element group 140:  members (11) 
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_0/$entry
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_0/rr
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_3/rr
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_2/rr
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/$entry
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_3/$entry
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_2/$entry
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_1/$entry
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_1/rr
      -- CP-element group 140: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_sample_start_
      -- 
    rr_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(140), ack => ptr_deref_489_load_0_req_0); -- 
    rr_1802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(140), ack => ptr_deref_489_load_1_req_0); -- 
    rr_1807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(140), ack => ptr_deref_489_load_2_req_0); -- 
    rr_1812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(140), ack => ptr_deref_489_load_3_req_0); -- 
    testConfigure_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(142) & testConfigure_CP_684_elements(284);
      gj_testConfigure_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	145 
    -- CP-element group 141: 	147 
    -- CP-element group 141: 	149 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	208 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_sample_complete
      -- 
    testConfigure_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(143) & testConfigure_CP_684_elements(145) & testConfigure_CP_684_elements(147) & testConfigure_CP_684_elements(149);
      gj_testConfigure_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  transition  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: 	146 
    -- CP-element group 142: 	148 
    -- CP-element group 142: 	150 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_update_complete
      -- 
    testConfigure_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(144) & testConfigure_CP_684_elements(146) & testConfigure_CP_684_elements(148) & testConfigure_CP_684_elements(150);
      gj_testConfigure_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	284 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_0_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_0_Sample/$exit
      -- 
    ra_1752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_addr_0_ack_0, ack => testConfigure_CP_684_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	284 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	142 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_0_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_0_Update/$exit
      -- 
    ca_1757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_addr_0_ack_1, ack => testConfigure_CP_684_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	284 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	141 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_1_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_1_Sample/$exit
      -- 
    ra_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_addr_1_ack_0, ack => testConfigure_CP_684_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	284 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	142 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_1_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_1_Update/$exit
      -- 
    ca_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_addr_1_ack_1, ack => testConfigure_CP_684_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	284 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	141 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_2_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_2_Sample/$exit
      -- 
    ra_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_addr_2_ack_0, ack => testConfigure_CP_684_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	284 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	142 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_2_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_2_Update/$exit
      -- 
    ca_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_addr_2_ack_1, ack => testConfigure_CP_684_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	284 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	141 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_3_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_3_Sample/$exit
      -- 
    ra_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_addr_3_ack_0, ack => testConfigure_CP_684_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	284 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	142 
    -- CP-element group 150:  members (2) 
      -- CP-element group 150: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_3_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_3_Update/$exit
      -- 
    ca_1787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_addr_3_ack_1, ack => testConfigure_CP_684_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	140 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	155 
    -- CP-element group 151:  members (2) 
      -- CP-element group 151: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_0/$exit
      -- CP-element group 151: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_0/ra
      -- 
    ra_1798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_load_0_ack_0, ack => testConfigure_CP_684_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	140 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_1/ra
      -- CP-element group 152: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_1/$exit
      -- 
    ra_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_load_1_ack_0, ack => testConfigure_CP_684_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	140 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_2/$exit
      -- CP-element group 153: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_2/ra
      -- 
    ra_1808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_load_2_ack_0, ack => testConfigure_CP_684_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	140 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (2) 
      -- CP-element group 154: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_3/$exit
      -- CP-element group 154: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/word_3/ra
      -- 
    ra_1813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_load_3_ack_0, ack => testConfigure_CP_684_elements(154)); -- 
    -- CP-element group 155:  join  transition  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	151 
    -- CP-element group 155: 	152 
    -- CP-element group 155: 	153 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Sample/word_access_start/$exit
      -- CP-element group 155: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_sample_completed_
      -- 
    testConfigure_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(151) & testConfigure_CP_684_elements(152) & testConfigure_CP_684_elements(153) & testConfigure_CP_684_elements(154);
      gj_testConfigure_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	284 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	160 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_0/$exit
      -- CP-element group 156: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_0/ca
      -- 
    ca_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_load_0_ack_1, ack => testConfigure_CP_684_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	284 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	160 
    -- CP-element group 157:  members (2) 
      -- CP-element group 157: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_1/$exit
      -- CP-element group 157: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_1/ca
      -- 
    ca_1829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_load_1_ack_1, ack => testConfigure_CP_684_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	284 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (2) 
      -- CP-element group 158: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_2/$exit
      -- CP-element group 158: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_2/ca
      -- 
    ca_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_load_2_ack_1, ack => testConfigure_CP_684_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	284 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_3/$exit
      -- CP-element group 159: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_3/ca
      -- 
    ca_1839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_489_load_3_ack_1, ack => testConfigure_CP_684_elements(159)); -- 
    -- CP-element group 160:  join  transition  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	156 
    -- CP-element group 160: 	157 
    -- CP-element group 160: 	158 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	203 
    -- CP-element group 160:  members (7) 
      -- CP-element group 160: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/$exit
      -- CP-element group 160: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/ptr_deref_489_Merge/$entry
      -- CP-element group 160: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/ptr_deref_489_Merge/$exit
      -- CP-element group 160: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/ptr_deref_489_Merge/merge_req
      -- CP-element group 160: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/ptr_deref_489_Merge/merge_ack
      -- 
    testConfigure_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(156) & testConfigure_CP_684_elements(157) & testConfigure_CP_684_elements(158) & testConfigure_CP_684_elements(159);
      gj_testConfigure_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  fork  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	284 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	172 
    -- CP-element group 161: 	173 
    -- CP-element group 161: 	174 
    -- CP-element group 161: 	175 
    -- CP-element group 161:  members (11) 
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_2/$entry
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_2/rr
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_3/$entry
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_3/rr
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_1/rr
      -- CP-element group 161: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_1/$entry
      -- 
    rr_1916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(161), ack => ptr_deref_501_load_0_req_0); -- 
    rr_1921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(161), ack => ptr_deref_501_load_1_req_0); -- 
    rr_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(161), ack => ptr_deref_501_load_2_req_0); -- 
    rr_1931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(161), ack => ptr_deref_501_load_3_req_0); -- 
    testConfigure_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(163) & testConfigure_CP_684_elements(284);
      gj_testConfigure_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  join  transition  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: 	166 
    -- CP-element group 162: 	168 
    -- CP-element group 162: 	170 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	208 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_sample_complete
      -- 
    testConfigure_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(164) & testConfigure_CP_684_elements(166) & testConfigure_CP_684_elements(168) & testConfigure_CP_684_elements(170);
      gj_testConfigure_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: 	167 
    -- CP-element group 163: 	169 
    -- CP-element group 163: 	171 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_address_calculated
      -- CP-element group 163: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_update_complete
      -- 
    testConfigure_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(165) & testConfigure_CP_684_elements(167) & testConfigure_CP_684_elements(169) & testConfigure_CP_684_elements(171);
      gj_testConfigure_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	284 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_0_Sample/ra
      -- CP-element group 164: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_0_Sample/$exit
      -- 
    ra_1871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_addr_0_ack_0, ack => testConfigure_CP_684_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	284 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_0_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_0_Update/$exit
      -- 
    ca_1876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_addr_0_ack_1, ack => testConfigure_CP_684_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	284 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	162 
    -- CP-element group 166:  members (2) 
      -- CP-element group 166: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_1_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_1_Sample/$exit
      -- 
    ra_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_addr_1_ack_0, ack => testConfigure_CP_684_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	284 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	163 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_1_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_1_Update/$exit
      -- 
    ca_1886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_addr_1_ack_1, ack => testConfigure_CP_684_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	284 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	162 
    -- CP-element group 168:  members (2) 
      -- CP-element group 168: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_2_Sample/ra
      -- CP-element group 168: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_2_Sample/$exit
      -- 
    ra_1891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_addr_2_ack_0, ack => testConfigure_CP_684_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	284 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	163 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_2_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_2_Update/$exit
      -- 
    ca_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_addr_2_ack_1, ack => testConfigure_CP_684_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	284 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	162 
    -- CP-element group 170:  members (2) 
      -- CP-element group 170: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_3_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_3_Sample/$exit
      -- 
    ra_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_addr_3_ack_0, ack => testConfigure_CP_684_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	284 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	163 
    -- CP-element group 171:  members (2) 
      -- CP-element group 171: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_3_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_3_Update/$exit
      -- 
    ca_1906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_addr_3_ack_1, ack => testConfigure_CP_684_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	161 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	176 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_0/$exit
      -- CP-element group 172: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_0/ra
      -- 
    ra_1917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_0_ack_0, ack => testConfigure_CP_684_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	161 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	176 
    -- CP-element group 173:  members (2) 
      -- CP-element group 173: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_1/ra
      -- CP-element group 173: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_1/$exit
      -- 
    ra_1922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_1_ack_0, ack => testConfigure_CP_684_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	161 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (2) 
      -- CP-element group 174: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_2/$exit
      -- CP-element group 174: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_2/ra
      -- 
    ra_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_2_ack_0, ack => testConfigure_CP_684_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	161 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (2) 
      -- CP-element group 175: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_3/$exit
      -- CP-element group 175: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/word_3/ra
      -- 
    ra_1932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_3_ack_0, ack => testConfigure_CP_684_elements(175)); -- 
    -- CP-element group 176:  join  transition  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	172 
    -- CP-element group 176: 	173 
    -- CP-element group 176: 	174 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/word_access_start/$exit
      -- CP-element group 176: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_sample_completed_
      -- 
    testConfigure_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(172) & testConfigure_CP_684_elements(173) & testConfigure_CP_684_elements(174) & testConfigure_CP_684_elements(175);
      gj_testConfigure_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	284 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	181 
    -- CP-element group 177:  members (2) 
      -- CP-element group 177: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_0/ca
      -- CP-element group 177: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_0/$exit
      -- 
    ca_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_0_ack_1, ack => testConfigure_CP_684_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	284 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_1/$exit
      -- CP-element group 178: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_1/ca
      -- 
    ca_1948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_1_ack_1, ack => testConfigure_CP_684_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	284 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_2/$exit
      -- CP-element group 179: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_2/ca
      -- 
    ca_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_2_ack_1, ack => testConfigure_CP_684_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	284 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_3/$exit
      -- CP-element group 180: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_3/ca
      -- 
    ca_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_501_load_3_ack_1, ack => testConfigure_CP_684_elements(180)); -- 
    -- CP-element group 181:  join  transition  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	177 
    -- CP-element group 181: 	178 
    -- CP-element group 181: 	179 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	203 
    -- CP-element group 181:  members (7) 
      -- CP-element group 181: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/ptr_deref_501_Merge/merge_ack
      -- CP-element group 181: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/$exit
      -- CP-element group 181: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/ptr_deref_501_Merge/merge_req
      -- CP-element group 181: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/ptr_deref_501_Merge/$exit
      -- CP-element group 181: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/ptr_deref_501_Merge/$entry
      -- 
    testConfigure_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(177) & testConfigure_CP_684_elements(178) & testConfigure_CP_684_elements(179) & testConfigure_CP_684_elements(180);
      gj_testConfigure_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  fork  transition  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	284 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	193 
    -- CP-element group 182: 	194 
    -- CP-element group 182: 	195 
    -- CP-element group 182: 	196 
    -- CP-element group 182:  members (11) 
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_0/rr
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_3/rr
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_1/rr
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_2/$entry
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_2/rr
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_3/$entry
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/$entry
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_0/$entry
      -- CP-element group 182: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_1/$entry
      -- 
    rr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(182), ack => ptr_deref_513_load_0_req_0); -- 
    rr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(182), ack => ptr_deref_513_load_1_req_0); -- 
    rr_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(182), ack => ptr_deref_513_load_2_req_0); -- 
    rr_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(182), ack => ptr_deref_513_load_3_req_0); -- 
    testConfigure_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(184) & testConfigure_CP_684_elements(284);
      gj_testConfigure_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: 	187 
    -- CP-element group 183: 	189 
    -- CP-element group 183: 	191 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	208 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_sample_complete
      -- 
    testConfigure_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(185) & testConfigure_CP_684_elements(187) & testConfigure_CP_684_elements(189) & testConfigure_CP_684_elements(191);
      gj_testConfigure_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  join  transition  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: 	188 
    -- CP-element group 184: 	190 
    -- CP-element group 184: 	192 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (2) 
      -- CP-element group 184: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_update_complete
      -- CP-element group 184: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_address_calculated
      -- 
    testConfigure_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(186) & testConfigure_CP_684_elements(188) & testConfigure_CP_684_elements(190) & testConfigure_CP_684_elements(192);
      gj_testConfigure_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	284 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	183 
    -- CP-element group 185:  members (2) 
      -- CP-element group 185: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_0_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_0_Sample/$exit
      -- 
    ra_1990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_addr_0_ack_0, ack => testConfigure_CP_684_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	284 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (2) 
      -- CP-element group 186: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_0_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_0_Update/ca
      -- 
    ca_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_addr_0_ack_1, ack => testConfigure_CP_684_elements(186)); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	284 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	183 
    -- CP-element group 187:  members (2) 
      -- CP-element group 187: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_1_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_1_Sample/$exit
      -- 
    ra_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_addr_1_ack_0, ack => testConfigure_CP_684_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	284 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	184 
    -- CP-element group 188:  members (2) 
      -- CP-element group 188: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_1_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_1_Update/ca
      -- 
    ca_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_addr_1_ack_1, ack => testConfigure_CP_684_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	284 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	183 
    -- CP-element group 189:  members (2) 
      -- CP-element group 189: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_2_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_2_Sample/$exit
      -- 
    ra_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_addr_2_ack_0, ack => testConfigure_CP_684_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	284 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	184 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_2_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_2_Update/ca
      -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_addr_2_ack_1, ack => testConfigure_CP_684_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	284 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	183 
    -- CP-element group 191:  members (2) 
      -- CP-element group 191: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_3_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_3_Sample/ra
      -- 
    ra_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_addr_3_ack_0, ack => testConfigure_CP_684_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	284 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	184 
    -- CP-element group 192:  members (2) 
      -- CP-element group 192: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_3_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_3_Update/$exit
      -- 
    ca_2025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_addr_3_ack_1, ack => testConfigure_CP_684_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	182 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	197 
    -- CP-element group 193:  members (2) 
      -- CP-element group 193: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_0/ra
      -- CP-element group 193: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_0/$exit
      -- 
    ra_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_0_ack_0, ack => testConfigure_CP_684_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	182 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (2) 
      -- CP-element group 194: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_1/$exit
      -- CP-element group 194: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_1/ra
      -- 
    ra_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_1_ack_0, ack => testConfigure_CP_684_elements(194)); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	182 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (2) 
      -- CP-element group 195: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_2/$exit
      -- CP-element group 195: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_2/ra
      -- 
    ra_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_2_ack_0, ack => testConfigure_CP_684_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	182 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (2) 
      -- CP-element group 196: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_3/$exit
      -- CP-element group 196: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/word_3/ra
      -- 
    ra_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_3_ack_0, ack => testConfigure_CP_684_elements(196)); -- 
    -- CP-element group 197:  join  transition  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	193 
    -- CP-element group 197: 	194 
    -- CP-element group 197: 	195 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/word_access_start/$exit
      -- CP-element group 197: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Sample/$exit
      -- 
    testConfigure_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(193) & testConfigure_CP_684_elements(194) & testConfigure_CP_684_elements(195) & testConfigure_CP_684_elements(196);
      gj_testConfigure_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	284 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	202 
    -- CP-element group 198:  members (2) 
      -- CP-element group 198: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_0/$exit
      -- CP-element group 198: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_0/ca
      -- 
    ca_2062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_0_ack_1, ack => testConfigure_CP_684_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	284 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	202 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_1/$exit
      -- CP-element group 199: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_1/ca
      -- 
    ca_2067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_1_ack_1, ack => testConfigure_CP_684_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	284 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (2) 
      -- CP-element group 200: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_2/$exit
      -- CP-element group 200: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_2/ca
      -- 
    ca_2072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_2_ack_1, ack => testConfigure_CP_684_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	284 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (2) 
      -- CP-element group 201: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_3/$exit
      -- CP-element group 201: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_3/ca
      -- 
    ca_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_513_load_3_ack_1, ack => testConfigure_CP_684_elements(201)); -- 
    -- CP-element group 202:  join  transition  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	198 
    -- CP-element group 202: 	199 
    -- CP-element group 202: 	200 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (7) 
      -- CP-element group 202: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/$exit
      -- CP-element group 202: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/ptr_deref_513_Merge/$entry
      -- CP-element group 202: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/ptr_deref_513_Merge/$exit
      -- CP-element group 202: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/ptr_deref_513_Merge/merge_req
      -- CP-element group 202: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/ptr_deref_513_Merge/merge_ack
      -- 
    testConfigure_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(198) & testConfigure_CP_684_elements(199) & testConfigure_CP_684_elements(200) & testConfigure_CP_684_elements(201);
      gj_testConfigure_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	160 
    -- CP-element group 203: 	181 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_Sample/rr
      -- 
    rr_2090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(203), ack => type_cast_527_inst_req_0); -- 
    testConfigure_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(160) & testConfigure_CP_684_elements(181) & testConfigure_CP_684_elements(202);
      gj_testConfigure_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_Sample/ra
      -- 
    ra_2091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_527_inst_ack_0, ack => testConfigure_CP_684_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	284 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	208 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_Update/ca
      -- 
    ca_2096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_527_inst_ack_1, ack => testConfigure_CP_684_elements(205)); -- 
    -- CP-element group 206:  transition  delay-element  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	124 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	130 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_ptr_deref_457_delay
      -- 
    -- Element group testConfigure_CP_684_elements(206) is a control-delay.
    cp_element_206_delay: control_delay_element  generic map(name => " 206_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(124), ack => testConfigure_CP_684_elements(206), clk => clk, reset =>reset);
    -- CP-element group 207:  transition  delay-element  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	131 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	137 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_ptr_deref_476_delay
      -- 
    -- Element group testConfigure_CP_684_elements(207) is a control-delay.
    cp_element_207_delay: control_delay_element  generic map(name => " 207_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(131), ack => testConfigure_CP_684_elements(207), clk => clk, reset =>reset);
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	118 
    -- CP-element group 208: 	125 
    -- CP-element group 208: 	132 
    -- CP-element group 208: 	139 
    -- CP-element group 208: 	141 
    -- CP-element group 208: 	162 
    -- CP-element group 208: 	183 
    -- CP-element group 208: 	205 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_275/if_stmt_541__entry__
      -- CP-element group 208: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540__exit__
      -- CP-element group 208: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/$exit
      -- CP-element group 208: 	 branch_block_stmt_275/if_stmt_541_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_275/if_stmt_541_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_275/if_stmt_541_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_275/if_stmt_541_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_275/R_cmp2583_542_place
      -- CP-element group 208: 	 branch_block_stmt_275/if_stmt_541_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_275/if_stmt_541_else_link/$entry
      -- 
    branch_req_2106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(208), ack => if_stmt_541_branch_req_0); -- 
    testConfigure_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(118) & testConfigure_CP_684_elements(125) & testConfigure_CP_684_elements(132) & testConfigure_CP_684_elements(139) & testConfigure_CP_684_elements(141) & testConfigure_CP_684_elements(162) & testConfigure_CP_684_elements(183) & testConfigure_CP_684_elements(205);
      gj_testConfigure_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	291 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_275/if_stmt_541_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_275/if_stmt_541_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_275/forx_xend_forx_xend78
      -- CP-element group 209: 	 branch_block_stmt_275/forx_xend_forx_xend78_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_275/forx_xend_forx_xend78_PhiReq/$exit
      -- 
    if_choice_transition_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_541_branch_ack_1, ack => testConfigure_CP_684_elements(209)); -- 
    -- CP-element group 210:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (18) 
      -- CP-element group 210: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580__entry__
      -- CP-element group 210: 	 branch_block_stmt_275/merge_stmt_547__exit__
      -- CP-element group 210: 	 branch_block_stmt_275/if_stmt_541_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_275/if_stmt_541_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_275/forx_xend_bbx_xnph
      -- CP-element group 210: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/$entry
      -- CP-element group 210: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_update_start_
      -- CP-element group 210: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_Update/cr
      -- CP-element group 210: 	 branch_block_stmt_275/forx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_275/forx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_275/merge_stmt_547_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_275/merge_stmt_547_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_275/merge_stmt_547_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_275/merge_stmt_547_PhiAck/dummy
      -- 
    else_choice_transition_2115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_541_branch_ack_0, ack => testConfigure_CP_684_elements(210)); -- 
    rr_2128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(210), ack => type_cast_560_inst_req_0); -- 
    cr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(210), ack => type_cast_560_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_Sample/ra
      -- 
    ra_2129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_560_inst_ack_0, ack => testConfigure_CP_684_elements(211)); -- 
    -- CP-element group 212:  transition  place  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	285 
    -- CP-element group 212:  members (9) 
      -- CP-element group 212: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27
      -- CP-element group 212: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580__exit__
      -- CP-element group 212: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/$exit
      -- CP-element group 212: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_275/assign_stmt_552_to_assign_stmt_580/type_cast_560_Update/ca
      -- CP-element group 212: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27_PhiReq/phi_stmt_583/$entry
      -- CP-element group 212: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/$entry
      -- 
    ca_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_560_inst_ack_1, ack => testConfigure_CP_684_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	290 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	252 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_sample_complete
      -- CP-element group 213: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_Sample/ack
      -- 
    ack_2163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_595_index_offset_ack_0, ack => testConfigure_CP_684_elements(213)); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	290 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (11) 
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_root_address_calculated
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_offset_calculated
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_Update/ack
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_base_plus_offset/$entry
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_base_plus_offset/$exit
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_base_plus_offset/sum_rename_req
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_base_plus_offset/sum_rename_ack
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_request/$entry
      -- CP-element group 214: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_request/req
      -- 
    ack_2168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_595_index_offset_ack_1, ack => testConfigure_CP_684_elements(214)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(214), ack => addr_of_596_final_reg_req_0); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_request/$exit
      -- CP-element group 215: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_request/ack
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_596_final_reg_ack_0, ack => testConfigure_CP_684_elements(215)); -- 
    -- CP-element group 216:  fork  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	290 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	249 
    -- CP-element group 216:  members (19) 
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_complete/$exit
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_complete/ack
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_address_calculated
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_word_address_calculated
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_root_address_calculated
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_address_resized
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_addr_resize/$entry
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_addr_resize/$exit
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_addr_resize/base_resize_req
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_addr_resize/base_resize_ack
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_plus_offset/$entry
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_plus_offset/$exit
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_plus_offset/sum_rename_req
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_base_plus_offset/sum_rename_ack
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_word_addrgen/$entry
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_word_addrgen/$exit
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_word_addrgen/root_register_req
      -- CP-element group 216: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_word_addrgen/root_register_ack
      -- 
    ack_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_596_final_reg_ack_1, ack => testConfigure_CP_684_elements(216)); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	290 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_update_start_
      -- CP-element group 217: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_Update/cr
      -- 
    ra_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_599_inst_ack_0, ack => testConfigure_CP_684_elements(217)); -- 
    cr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(217), ack => RPIPE_zeropad_input_pipe_599_inst_req_1); -- 
    -- CP-element group 218:  fork  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (9) 
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_Sample/rr
      -- 
    ca_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_599_inst_ack_1, ack => testConfigure_CP_684_elements(218)); -- 
    rr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(218), ack => type_cast_603_inst_req_0); -- 
    rr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(218), ack => RPIPE_zeropad_input_pipe_612_inst_req_0); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_Sample/ra
      -- 
    ra_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_603_inst_ack_0, ack => testConfigure_CP_684_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	290 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	249 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_Update/ca
      -- 
    ca_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_603_inst_ack_1, ack => testConfigure_CP_684_elements(220)); -- 
    -- CP-element group 221:  transition  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (6) 
      -- CP-element group 221: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_update_start_
      -- CP-element group 221: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_Sample/ra
      -- CP-element group 221: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_Update/cr
      -- 
    ra_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_612_inst_ack_0, ack => testConfigure_CP_684_elements(221)); -- 
    cr_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(221), ack => RPIPE_zeropad_input_pipe_612_inst_req_1); -- 
    -- CP-element group 222:  fork  transition  input  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222: 	225 
    -- CP-element group 222:  members (9) 
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_612_Update/ca
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_Sample/rr
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_Sample/rr
      -- 
    ca_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_612_inst_ack_1, ack => testConfigure_CP_684_elements(222)); -- 
    rr_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(222), ack => type_cast_616_inst_req_0); -- 
    rr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(222), ack => RPIPE_zeropad_input_pipe_630_inst_req_0); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_Sample/ra
      -- 
    ra_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_0, ack => testConfigure_CP_684_elements(223)); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	290 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	249 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_Update/ca
      -- 
    ca_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_1, ack => testConfigure_CP_684_elements(224)); -- 
    -- CP-element group 225:  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	222 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (6) 
      -- CP-element group 225: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_update_start_
      -- CP-element group 225: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_Sample/ra
      -- CP-element group 225: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_Update/cr
      -- 
    ra_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_630_inst_ack_0, ack => testConfigure_CP_684_elements(225)); -- 
    cr_2252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(225), ack => RPIPE_zeropad_input_pipe_630_inst_req_1); -- 
    -- CP-element group 226:  fork  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226: 	229 
    -- CP-element group 226:  members (9) 
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_630_Update/ca
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_Sample/rr
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_Sample/rr
      -- 
    ca_2253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_630_inst_ack_1, ack => testConfigure_CP_684_elements(226)); -- 
    rr_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(226), ack => type_cast_634_inst_req_0); -- 
    rr_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(226), ack => RPIPE_zeropad_input_pipe_648_inst_req_0); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_Sample/ra
      -- 
    ra_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_634_inst_ack_0, ack => testConfigure_CP_684_elements(227)); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	290 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	249 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_Update/ca
      -- 
    ca_2267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_634_inst_ack_1, ack => testConfigure_CP_684_elements(228)); -- 
    -- CP-element group 229:  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	226 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (6) 
      -- CP-element group 229: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_sample_completed_
      -- CP-element group 229: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_update_start_
      -- CP-element group 229: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_Sample/ra
      -- CP-element group 229: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_Update/cr
      -- 
    ra_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_648_inst_ack_0, ack => testConfigure_CP_684_elements(229)); -- 
    cr_2280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(229), ack => RPIPE_zeropad_input_pipe_648_inst_req_1); -- 
    -- CP-element group 230:  fork  transition  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230: 	233 
    -- CP-element group 230:  members (9) 
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_648_Update/ca
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_Sample/rr
      -- 
    ca_2281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_648_inst_ack_1, ack => testConfigure_CP_684_elements(230)); -- 
    rr_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(230), ack => type_cast_652_inst_req_0); -- 
    rr_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(230), ack => RPIPE_zeropad_input_pipe_666_inst_req_0); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_Sample/ra
      -- 
    ra_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_0, ack => testConfigure_CP_684_elements(231)); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	290 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	249 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_Update/ca
      -- 
    ca_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_1, ack => testConfigure_CP_684_elements(232)); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	230 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_update_start_
      -- CP-element group 233: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_Sample/ra
      -- CP-element group 233: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_Update/cr
      -- 
    ra_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_666_inst_ack_0, ack => testConfigure_CP_684_elements(233)); -- 
    cr_2308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(233), ack => RPIPE_zeropad_input_pipe_666_inst_req_1); -- 
    -- CP-element group 234:  fork  transition  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	237 
    -- CP-element group 234:  members (9) 
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_666_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_Sample/rr
      -- 
    ca_2309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_666_inst_ack_1, ack => testConfigure_CP_684_elements(234)); -- 
    rr_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(234), ack => type_cast_670_inst_req_0); -- 
    rr_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(234), ack => RPIPE_zeropad_input_pipe_684_inst_req_0); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_Sample/ra
      -- 
    ra_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_670_inst_ack_0, ack => testConfigure_CP_684_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	290 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	249 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_Update/ca
      -- 
    ca_2323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_670_inst_ack_1, ack => testConfigure_CP_684_elements(236)); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	234 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_update_start_
      -- CP-element group 237: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_Sample/ra
      -- CP-element group 237: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_Update/cr
      -- 
    ra_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_684_inst_ack_0, ack => testConfigure_CP_684_elements(237)); -- 
    cr_2336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(237), ack => RPIPE_zeropad_input_pipe_684_inst_req_1); -- 
    -- CP-element group 238:  fork  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: 	241 
    -- CP-element group 238:  members (9) 
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_684_Update/ca
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_Sample/rr
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_Sample/rr
      -- 
    ca_2337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_684_inst_ack_1, ack => testConfigure_CP_684_elements(238)); -- 
    rr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(238), ack => type_cast_688_inst_req_0); -- 
    rr_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(238), ack => RPIPE_zeropad_input_pipe_702_inst_req_0); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_Sample/ra
      -- 
    ra_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_0, ack => testConfigure_CP_684_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	290 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	249 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_Update/ca
      -- 
    ca_2351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_1, ack => testConfigure_CP_684_elements(240)); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	238 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_update_start_
      -- CP-element group 241: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_Sample/ra
      -- CP-element group 241: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_Update/cr
      -- 
    ra_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_702_inst_ack_0, ack => testConfigure_CP_684_elements(241)); -- 
    cr_2364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(241), ack => RPIPE_zeropad_input_pipe_702_inst_req_1); -- 
    -- CP-element group 242:  fork  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242: 	245 
    -- CP-element group 242:  members (9) 
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_702_Update/ca
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_Sample/rr
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_Sample/rr
      -- 
    ca_2365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_702_inst_ack_1, ack => testConfigure_CP_684_elements(242)); -- 
    rr_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(242), ack => type_cast_706_inst_req_0); -- 
    rr_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(242), ack => RPIPE_zeropad_input_pipe_720_inst_req_0); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_Sample/ra
      -- 
    ra_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_706_inst_ack_0, ack => testConfigure_CP_684_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	290 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	249 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_Update/ca
      -- 
    ca_2379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_706_inst_ack_1, ack => testConfigure_CP_684_elements(244)); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	242 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_update_start_
      -- CP-element group 245: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_Sample/ra
      -- CP-element group 245: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_Update/cr
      -- 
    ra_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_720_inst_ack_0, ack => testConfigure_CP_684_elements(245)); -- 
    cr_2392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(245), ack => RPIPE_zeropad_input_pipe_720_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_720_Update/ca
      -- CP-element group 246: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_Sample/rr
      -- 
    ca_2393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_720_inst_ack_1, ack => testConfigure_CP_684_elements(246)); -- 
    rr_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(246), ack => type_cast_724_inst_req_0); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_Sample/ra
      -- 
    ra_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_724_inst_ack_0, ack => testConfigure_CP_684_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	290 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_Update/ca
      -- 
    ca_2407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_724_inst_ack_1, ack => testConfigure_CP_684_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	216 
    -- CP-element group 249: 	220 
    -- CP-element group 249: 	224 
    -- CP-element group 249: 	228 
    -- CP-element group 249: 	232 
    -- CP-element group 249: 	236 
    -- CP-element group 249: 	240 
    -- CP-element group 249: 	244 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (9) 
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/ptr_deref_732_Split/$entry
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/ptr_deref_732_Split/$exit
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/ptr_deref_732_Split/split_req
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/ptr_deref_732_Split/split_ack
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/word_access_start/$entry
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/word_access_start/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/word_access_start/word_0/rr
      -- 
    rr_2445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(249), ack => ptr_deref_732_store_0_req_0); -- 
    testConfigure_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(216) & testConfigure_CP_684_elements(220) & testConfigure_CP_684_elements(224) & testConfigure_CP_684_elements(228) & testConfigure_CP_684_elements(232) & testConfigure_CP_684_elements(236) & testConfigure_CP_684_elements(240) & testConfigure_CP_684_elements(244) & testConfigure_CP_684_elements(248);
      gj_testConfigure_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (5) 
      -- CP-element group 250: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/word_access_start/$exit
      -- CP-element group 250: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/word_access_start/word_0/$exit
      -- CP-element group 250: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Sample/word_access_start/word_0/ra
      -- 
    ra_2446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_732_store_0_ack_0, ack => testConfigure_CP_684_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	290 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (5) 
      -- CP-element group 251: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Update/word_access_complete/$exit
      -- CP-element group 251: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Update/word_access_complete/word_0/$exit
      -- CP-element group 251: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Update/word_access_complete/word_0/ca
      -- 
    ca_2457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_732_store_0_ack_1, ack => testConfigure_CP_684_elements(251)); -- 
    -- CP-element group 252:  branch  join  transition  place  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	213 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (10) 
      -- CP-element group 252: 	 branch_block_stmt_275/if_stmt_746__entry__
      -- CP-element group 252: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745__exit__
      -- CP-element group 252: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/$exit
      -- CP-element group 252: 	 branch_block_stmt_275/if_stmt_746_dead_link/$entry
      -- CP-element group 252: 	 branch_block_stmt_275/if_stmt_746_eval_test/$entry
      -- CP-element group 252: 	 branch_block_stmt_275/if_stmt_746_eval_test/$exit
      -- CP-element group 252: 	 branch_block_stmt_275/if_stmt_746_eval_test/branch_req
      -- CP-element group 252: 	 branch_block_stmt_275/R_exitcond10_747_place
      -- CP-element group 252: 	 branch_block_stmt_275/if_stmt_746_if_link/$entry
      -- CP-element group 252: 	 branch_block_stmt_275/if_stmt_746_else_link/$entry
      -- 
    branch_req_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(252), ack => if_stmt_746_branch_req_0); -- 
    testConfigure_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(213) & testConfigure_CP_684_elements(251);
      gj_testConfigure_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  merge  transition  place  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	291 
    -- CP-element group 253:  members (13) 
      -- CP-element group 253: 	 branch_block_stmt_275/forx_xend78x_xloopexit_forx_xend78
      -- CP-element group 253: 	 branch_block_stmt_275/merge_stmt_752__exit__
      -- CP-element group 253: 	 branch_block_stmt_275/if_stmt_746_if_link/$exit
      -- CP-element group 253: 	 branch_block_stmt_275/if_stmt_746_if_link/if_choice_transition
      -- CP-element group 253: 	 branch_block_stmt_275/forx_xbody27_forx_xend78x_xloopexit
      -- CP-element group 253: 	 branch_block_stmt_275/forx_xbody27_forx_xend78x_xloopexit_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_275/forx_xbody27_forx_xend78x_xloopexit_PhiReq/$exit
      -- CP-element group 253: 	 branch_block_stmt_275/merge_stmt_752_PhiReqMerge
      -- CP-element group 253: 	 branch_block_stmt_275/merge_stmt_752_PhiAck/$entry
      -- CP-element group 253: 	 branch_block_stmt_275/merge_stmt_752_PhiAck/$exit
      -- CP-element group 253: 	 branch_block_stmt_275/merge_stmt_752_PhiAck/dummy
      -- CP-element group 253: 	 branch_block_stmt_275/forx_xend78x_xloopexit_forx_xend78_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_275/forx_xend78x_xloopexit_forx_xend78_PhiReq/$exit
      -- 
    if_choice_transition_2470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_746_branch_ack_1, ack => testConfigure_CP_684_elements(253)); -- 
    -- CP-element group 254:  fork  transition  place  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	286 
    -- CP-element group 254: 	287 
    -- CP-element group 254:  members (12) 
      -- CP-element group 254: 	 branch_block_stmt_275/if_stmt_746_else_link/$exit
      -- CP-element group 254: 	 branch_block_stmt_275/if_stmt_746_else_link/else_choice_transition
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/$entry
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/$entry
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/$entry
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/$entry
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/$entry
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/Sample/rr
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_746_branch_ack_0, ack => testConfigure_CP_684_elements(254)); -- 
    rr_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(254), ack => type_cast_589_inst_req_0); -- 
    cr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(254), ack => type_cast_589_inst_req_1); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	291 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_Sample/ra
      -- 
    ra_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_757_inst_ack_0, ack => testConfigure_CP_684_elements(255)); -- 
    -- CP-element group 256:  transition  place  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	291 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (16) 
      -- CP-element group 256: 	 branch_block_stmt_275/merge_stmt_760__exit__
      -- CP-element group 256: 	 branch_block_stmt_275/branch_block_stmt_275__exit__
      -- CP-element group 256: 	 branch_block_stmt_275/return__
      -- CP-element group 256: 	 branch_block_stmt_275/assign_stmt_758__exit__
      -- CP-element group 256: 	 branch_block_stmt_275/$exit
      -- CP-element group 256: 	 $exit
      -- CP-element group 256: 	 branch_block_stmt_275/return___PhiReq/$entry
      -- CP-element group 256: 	 branch_block_stmt_275/return___PhiReq/$exit
      -- CP-element group 256: 	 branch_block_stmt_275/merge_stmt_760_PhiAck/$entry
      -- CP-element group 256: 	 branch_block_stmt_275/merge_stmt_760_PhiAck/dummy
      -- CP-element group 256: 	 branch_block_stmt_275/merge_stmt_760_PhiAck/$exit
      -- CP-element group 256: 	 branch_block_stmt_275/merge_stmt_760_PhiReqMerge
      -- CP-element group 256: 	 branch_block_stmt_275/assign_stmt_758/$exit
      -- CP-element group 256: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_Update/ca
      -- 
    ca_2493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_757_inst_ack_1, ack => testConfigure_CP_684_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	115 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (2) 
      -- CP-element group 257: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/Sample/ra
      -- 
    ra_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_338_inst_ack_0, ack => testConfigure_CP_684_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	115 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/Update/ca
      -- 
    ca_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_338_inst_ack_1, ack => testConfigure_CP_684_elements(258)); -- 
    -- CP-element group 259:  join  transition  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	263 
    -- CP-element group 259:  members (5) 
      -- CP-element group 259: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/$exit
      -- CP-element group 259: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/$exit
      -- CP-element group 259: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/$exit
      -- CP-element group 259: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/SplitProtocol/$exit
      -- CP-element group 259: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_req
      -- 
    phi_stmt_335_req_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_335_req_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(259), ack => phi_stmt_335_req_0); -- 
    testConfigure_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(257) & testConfigure_CP_684_elements(258);
      gj_testConfigure_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	115 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (2) 
      -- CP-element group 260: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/Sample/ra
      -- 
    ra_2548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_0, ack => testConfigure_CP_684_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	115 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (2) 
      -- CP-element group 261: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/Update/ca
      -- 
    ca_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_1, ack => testConfigure_CP_684_elements(261)); -- 
    -- CP-element group 262:  join  transition  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (5) 
      -- CP-element group 262: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/$exit
      -- CP-element group 262: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/$exit
      -- CP-element group 262: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/$exit
      -- CP-element group 262: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_345/SplitProtocol/$exit
      -- CP-element group 262: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_req
      -- 
    phi_stmt_342_req_2554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_342_req_2554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(262), ack => phi_stmt_342_req_0); -- 
    testConfigure_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(260) & testConfigure_CP_684_elements(261);
      gj_testConfigure_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  join  transition  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	259 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	269 
    -- CP-element group 263:  members (1) 
      -- CP-element group 263: 	 branch_block_stmt_275/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(259) & testConfigure_CP_684_elements(262);
      gj_testConfigure_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  transition  output  delay-element  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	58 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	268 
    -- CP-element group 264:  members (4) 
      -- CP-element group 264: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_335/$exit
      -- CP-element group 264: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/$exit
      -- CP-element group 264: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_341_konst_delay_trans
      -- CP-element group 264: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_335/phi_stmt_335_req
      -- 
    phi_stmt_335_req_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_335_req_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(264), ack => phi_stmt_335_req_1); -- 
    -- Element group testConfigure_CP_684_elements(264) is a control-delay.
    cp_element_264_delay: control_delay_element  generic map(name => " 264_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(58), ack => testConfigure_CP_684_elements(264), clk => clk, reset =>reset);
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	58 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (2) 
      -- CP-element group 265: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/Sample/ra
      -- 
    ra_2582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_347_inst_ack_0, ack => testConfigure_CP_684_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	58 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/Update/ca
      -- 
    ca_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_347_inst_ack_1, ack => testConfigure_CP_684_elements(266)); -- 
    -- CP-element group 267:  join  transition  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (5) 
      -- CP-element group 267: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/$exit
      -- CP-element group 267: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/$exit
      -- CP-element group 267: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/$exit
      -- CP-element group 267: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_sources/type_cast_347/SplitProtocol/$exit
      -- CP-element group 267: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_342/phi_stmt_342_req
      -- 
    phi_stmt_342_req_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_342_req_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(267), ack => phi_stmt_342_req_1); -- 
    testConfigure_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(265) & testConfigure_CP_684_elements(266);
      gj_testConfigure_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  join  transition  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	264 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (1) 
      -- CP-element group 268: 	 branch_block_stmt_275/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(264) & testConfigure_CP_684_elements(267);
      gj_testConfigure_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  merge  fork  transition  place  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	263 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (2) 
      -- CP-element group 269: 	 branch_block_stmt_275/merge_stmt_334_PhiReqMerge
      -- CP-element group 269: 	 branch_block_stmt_275/merge_stmt_334_PhiAck/$entry
      -- 
    testConfigure_CP_684_elements(269) <= OrReduce(testConfigure_CP_684_elements(263) & testConfigure_CP_684_elements(268));
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (1) 
      -- CP-element group 270: 	 branch_block_stmt_275/merge_stmt_334_PhiAck/phi_stmt_335_ack
      -- 
    phi_stmt_335_ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_335_ack_0, ack => testConfigure_CP_684_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (1) 
      -- CP-element group 271: 	 branch_block_stmt_275/merge_stmt_334_PhiAck/phi_stmt_342_ack
      -- 
    phi_stmt_342_ack_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_342_ack_0, ack => testConfigure_CP_684_elements(271)); -- 
    -- CP-element group 272:  join  fork  transition  place  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	64 
    -- CP-element group 272: 	66 
    -- CP-element group 272: 	67 
    -- CP-element group 272: 	68 
    -- CP-element group 272: 	73 
    -- CP-element group 272: 	75 
    -- CP-element group 272: 	77 
    -- CP-element group 272: 	79 
    -- CP-element group 272: 	85 
    -- CP-element group 272: 	86 
    -- CP-element group 272: 	87 
    -- CP-element group 272: 	88 
    -- CP-element group 272: 	90 
    -- CP-element group 272: 	93 
    -- CP-element group 272: 	94 
    -- CP-element group 272: 	95 
    -- CP-element group 272: 	96 
    -- CP-element group 272: 	97 
    -- CP-element group 272: 	98 
    -- CP-element group 272: 	99 
    -- CP-element group 272: 	100 
    -- CP-element group 272: 	59 
    -- CP-element group 272: 	60 
    -- CP-element group 272: 	61 
    -- CP-element group 272: 	62 
    -- CP-element group 272: 	106 
    -- CP-element group 272: 	107 
    -- CP-element group 272: 	108 
    -- CP-element group 272: 	109 
    -- CP-element group 272: 	111 
    -- CP-element group 272:  members (97) 
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397__entry__
      -- CP-element group 272: 	 branch_block_stmt_275/merge_stmt_334__exit__
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_update_start_
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_357_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_update_start_
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_resized_1
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_computed_1
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_resize_1/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_resize_1/$exit
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_resize_1/index_resize_req
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_resize_1/index_resize_ack
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_sample_start
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_update_start
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_index_scale_1_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_update_start
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/array_obj_ref_363_final_index_sum_regn_Update/req
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_complete/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/addr_of_364_complete/req
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_update_start_
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/type_cast_368_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_update_start_
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_update_start
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_0_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_0_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_1_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_1_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_2_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_2_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_3_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_word_addrgen_3_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_0/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_0/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_1/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_1/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_2/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_2/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_3/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_371_Update/word_access_complete/word_3/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_update_start_
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_address_calculated
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_root_address_calculated
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_address_resized
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_addr_resize/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_addr_resize/$exit
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_addr_resize/base_resize_req
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_addr_resize/base_resize_ack
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_plus_offset/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_plus_offset/$exit
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_plus_offset/sum_rename_req
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_base_plus_offset/sum_rename_ack
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_sample_start
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_update_start
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_0_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_0_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_0_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_0_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_1_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_1_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_1_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_1_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_2_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_2_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_2_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_2_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_3_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_3_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_3_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_word_addrgen_3_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_0/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_0/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_1/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_1/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_2/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_2/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_3/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/ptr_deref_388_Update/word_access_complete/word_3/cr
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_275/assign_stmt_354_to_assign_stmt_397/RPIPE_zeropad_input_pipe_396_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_275/merge_stmt_334_PhiAck/$exit
      -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => type_cast_357_inst_req_0); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => type_cast_357_inst_req_1); -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => array_obj_ref_363_index_1_scale_req_0); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => array_obj_ref_363_index_1_scale_req_1); -- 
    req_1153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => array_obj_ref_363_index_offset_req_1); -- 
    req_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => addr_of_364_final_reg_req_1); -- 
    rr_1177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => type_cast_368_inst_req_0); -- 
    cr_1182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => type_cast_368_inst_req_1); -- 
    cr_1214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_371_addr_0_req_1); -- 
    cr_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_371_addr_1_req_1); -- 
    cr_1234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_371_addr_2_req_1); -- 
    cr_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_371_addr_3_req_1); -- 
    cr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_371_store_0_req_1); -- 
    cr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_371_store_1_req_1); -- 
    cr_1296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_371_store_2_req_1); -- 
    cr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_371_store_3_req_1); -- 
    rr_1328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_addr_0_req_0); -- 
    cr_1333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_addr_0_req_1); -- 
    rr_1338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_addr_1_req_0); -- 
    cr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_addr_1_req_1); -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_addr_2_req_0); -- 
    cr_1353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_addr_2_req_1); -- 
    rr_1358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_addr_3_req_0); -- 
    cr_1363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_addr_3_req_1); -- 
    cr_1400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_load_0_req_1); -- 
    cr_1405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_load_1_req_1); -- 
    cr_1410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_load_2_req_1); -- 
    cr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => ptr_deref_388_load_3_req_1); -- 
    rr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(272), ack => RPIPE_zeropad_input_pipe_396_inst_req_0); -- 
    testConfigure_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(270) & testConfigure_CP_684_elements(271);
      gj_testConfigure_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	116 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (2) 
      -- CP-element group 273: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/Sample/ra
      -- 
    ra_2618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_0, ack => testConfigure_CP_684_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	116 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/Update/ca
      -- 
    ca_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_1, ack => testConfigure_CP_684_elements(274)); -- 
    -- CP-element group 275:  join  transition  place  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (8) 
      -- CP-element group 275: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 275: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/$exit
      -- CP-element group 275: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/$exit
      -- CP-element group 275: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/$exit
      -- CP-element group 275: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_408/SplitProtocol/$exit
      -- CP-element group 275: 	 branch_block_stmt_275/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_405/phi_stmt_405_req
      -- CP-element group 275: 	 branch_block_stmt_275/merge_stmt_404_PhiReqMerge
      -- CP-element group 275: 	 branch_block_stmt_275/merge_stmt_404_PhiAck/$entry
      -- 
    phi_stmt_405_req_2624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_405_req_2624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(275), ack => phi_stmt_405_req_0); -- 
    testConfigure_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(273) & testConfigure_CP_684_elements(274);
      gj_testConfigure_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	280 
    -- CP-element group 276: 	281 
    -- CP-element group 276:  members (13) 
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend
      -- CP-element group 276: 	 branch_block_stmt_275/merge_stmt_404__exit__
      -- CP-element group 276: 	 branch_block_stmt_275/merge_stmt_404_PhiAck/$exit
      -- CP-element group 276: 	 branch_block_stmt_275/merge_stmt_404_PhiAck/phi_stmt_405_ack
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/$entry
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/$entry
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/$entry
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/$entry
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/Sample/rr
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/Update/$entry
      -- CP-element group 276: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/Update/cr
      -- 
    phi_stmt_405_ack_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_405_ack_0, ack => testConfigure_CP_684_elements(276)); -- 
    rr_2674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(276), ack => type_cast_417_inst_req_0); -- 
    cr_2679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(276), ack => type_cast_417_inst_req_1); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	57 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (2) 
      -- CP-element group 277: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/Sample/ra
      -- 
    ra_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_415_inst_ack_0, ack => testConfigure_CP_684_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	57 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/Update/ca
      -- 
    ca_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_415_inst_ack_1, ack => testConfigure_CP_684_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	283 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/$exit
      -- CP-element group 279: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/$exit
      -- CP-element group 279: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/$exit
      -- CP-element group 279: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/$exit
      -- CP-element group 279: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_415/SplitProtocol/$exit
      -- CP-element group 279: 	 branch_block_stmt_275/entry_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_req
      -- 
    phi_stmt_412_req_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_412_req_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(279), ack => phi_stmt_412_req_0); -- 
    testConfigure_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(277) & testConfigure_CP_684_elements(278);
      gj_testConfigure_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	276 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (2) 
      -- CP-element group 280: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/Sample/ra
      -- 
    ra_2675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_417_inst_ack_0, ack => testConfigure_CP_684_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	276 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/Update/ca
      -- 
    ca_2680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_417_inst_ack_1, ack => testConfigure_CP_684_elements(281)); -- 
    -- CP-element group 282:  join  transition  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (6) 
      -- CP-element group 282: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 282: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/$exit
      -- CP-element group 282: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/$exit
      -- CP-element group 282: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/$exit
      -- CP-element group 282: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_sources/type_cast_417/SplitProtocol/$exit
      -- CP-element group 282: 	 branch_block_stmt_275/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_412/phi_stmt_412_req
      -- 
    phi_stmt_412_req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_412_req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(282), ack => phi_stmt_412_req_1); -- 
    testConfigure_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(280) & testConfigure_CP_684_elements(281);
      gj_testConfigure_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  merge  transition  place  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	279 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (2) 
      -- CP-element group 283: 	 branch_block_stmt_275/merge_stmt_411_PhiReqMerge
      -- CP-element group 283: 	 branch_block_stmt_275/merge_stmt_411_PhiAck/$entry
      -- 
    testConfigure_CP_684_elements(283) <= OrReduce(testConfigure_CP_684_elements(279) & testConfigure_CP_684_elements(282));
    -- CP-element group 284:  fork  transition  place  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	117 
    -- CP-element group 284: 	118 
    -- CP-element group 284: 	119 
    -- CP-element group 284: 	122 
    -- CP-element group 284: 	123 
    -- CP-element group 284: 	125 
    -- CP-element group 284: 	129 
    -- CP-element group 284: 	130 
    -- CP-element group 284: 	132 
    -- CP-element group 284: 	136 
    -- CP-element group 284: 	137 
    -- CP-element group 284: 	139 
    -- CP-element group 284: 	140 
    -- CP-element group 284: 	143 
    -- CP-element group 284: 	144 
    -- CP-element group 284: 	145 
    -- CP-element group 284: 	146 
    -- CP-element group 284: 	147 
    -- CP-element group 284: 	148 
    -- CP-element group 284: 	149 
    -- CP-element group 284: 	150 
    -- CP-element group 284: 	156 
    -- CP-element group 284: 	157 
    -- CP-element group 284: 	158 
    -- CP-element group 284: 	159 
    -- CP-element group 284: 	161 
    -- CP-element group 284: 	164 
    -- CP-element group 284: 	165 
    -- CP-element group 284: 	166 
    -- CP-element group 284: 	167 
    -- CP-element group 284: 	168 
    -- CP-element group 284: 	169 
    -- CP-element group 284: 	170 
    -- CP-element group 284: 	171 
    -- CP-element group 284: 	177 
    -- CP-element group 284: 	178 
    -- CP-element group 284: 	179 
    -- CP-element group 284: 	180 
    -- CP-element group 284: 	182 
    -- CP-element group 284: 	185 
    -- CP-element group 284: 	186 
    -- CP-element group 284: 	187 
    -- CP-element group 284: 	188 
    -- CP-element group 284: 	189 
    -- CP-element group 284: 	190 
    -- CP-element group 284: 	191 
    -- CP-element group 284: 	192 
    -- CP-element group 284: 	198 
    -- CP-element group 284: 	199 
    -- CP-element group 284: 	200 
    -- CP-element group 284: 	201 
    -- CP-element group 284: 	205 
    -- CP-element group 284:  members (219) 
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_word_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_addr_resize/base_resize_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_addr_resize/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_addr_resize/base_resize_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_addr_resize/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_addr_resize/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_addr_resize/base_resize_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_addr_resize/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_word_addrgen/root_register_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540__entry__
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_addr_resize/base_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_275/merge_stmt_411__exit__
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_word_addrgen/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_addr_resize/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_word_addrgen/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_2/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_word_addrgen/root_register_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_address_resized
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_word_addrgen/root_register_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_addr_resize/base_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_word_addrgen/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_2_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_2_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_3/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_3/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_0_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_3_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_word_addrgen/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_addr_resize/base_resize_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_address_resized
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_1/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_addr_resize/base_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_address_resized
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_1/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_addr_resize/base_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_addr_resize/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_word_addrgen/root_register_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_sample_start
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_2/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_1/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_update_start
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_0_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_1/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_3_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_sample_start
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_1_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_1_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_2_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_2_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_3_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_3_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_1_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_1/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_1_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_2/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_2/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_0_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_3/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_Update/word_access_complete/word_3/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_address_resized
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_addr_resize/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_word_addrgen_0_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_update_start
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_3_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_3_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_3_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_3_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_base_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_3_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_476_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_word_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_2_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_addr_resize/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_3_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_addr_resize/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_3_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_3_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_base_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_2_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_2_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_2_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_2_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_2_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_2_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_1_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_address_resized
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_2_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_1_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_1_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_1_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_457_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_1_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_1_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_465_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_1_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_0_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_0_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_0_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_1_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_0_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_update_start
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_word_addrgen_sample_start
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_base_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_0_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_0_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_0_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_addr_resize/base_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_addr_resize/base_resize_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_489_base_addr_resize/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_501_word_addrgen_0_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_word_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/STORE_pad_419_Split/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/STORE_pad_419_Split/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/STORE_pad_419_Split/split_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/STORE_pad_419_Split/split_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/word_access_start/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/word_access_start/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Sample/word_access_start/word_0/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/STORE_pad_419_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/RPIPE_zeropad_input_pipe_423_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_427_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_word_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_address_resized
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_addr_resize/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_addr_resize/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_addr_resize/base_resize_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_addr_resize/base_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_word_addrgen/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_word_addrgen/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_word_addrgen/root_register_req
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_word_addrgen/root_register_ack
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_438_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_446_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_1/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_2/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_2/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_3/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/ptr_deref_513_Update/word_access_complete/word_3/cr
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_update_start_
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_275/assign_stmt_421_to_assign_stmt_540/type_cast_527_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_275/merge_stmt_411_PhiAck/$exit
      -- CP-element group 284: 	 branch_block_stmt_275/merge_stmt_411_PhiAck/phi_stmt_412_ack
      -- 
    phi_stmt_412_ack_2686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_412_ack_0, ack => testConfigure_CP_684_elements(284)); -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_addr_2_req_1); -- 
    cr_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_load_3_req_1); -- 
    cr_1947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_load_1_req_1); -- 
    cr_1724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_476_store_0_req_1); -- 
    cr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_load_0_req_1); -- 
    cr_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_load_2_req_1); -- 
    cr_1646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_457_store_0_req_1); -- 
    rr_1989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_addr_0_req_0); -- 
    cr_2024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_addr_3_req_1); -- 
    cr_2061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_load_0_req_1); -- 
    rr_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_addr_1_req_0); -- 
    rr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_addr_2_req_0); -- 
    rr_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_addr_3_req_0); -- 
    cr_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_addr_1_req_1); -- 
    cr_1828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_load_1_req_1); -- 
    cr_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_load_2_req_1); -- 
    cr_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_addr_0_req_1); -- 
    cr_1838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_load_3_req_1); -- 
    cr_1905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_addr_3_req_1); -- 
    cr_1786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_addr_3_req_1); -- 
    rr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_addr_3_req_0); -- 
    cr_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_addr_2_req_1); -- 
    rr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_addr_3_req_0); -- 
    cr_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_load_0_req_1); -- 
    cr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_addr_2_req_1); -- 
    rr_1890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_addr_2_req_0); -- 
    cr_1674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => type_cast_465_inst_req_1); -- 
    rr_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_addr_2_req_0); -- 
    cr_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_addr_1_req_1); -- 
    cr_1885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_addr_1_req_1); -- 
    rr_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_addr_1_req_0); -- 
    rr_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_addr_1_req_0); -- 
    cr_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_addr_0_req_1); -- 
    rr_1751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_489_addr_0_req_0); -- 
    cr_1875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_addr_0_req_1); -- 
    rr_1870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_501_addr_0_req_0); -- 
    rr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => STORE_pad_419_store_0_req_0); -- 
    cr_1490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => STORE_pad_419_store_0_req_1); -- 
    rr_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => RPIPE_zeropad_input_pipe_423_inst_req_0); -- 
    cr_1518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => type_cast_427_inst_req_1); -- 
    cr_1568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_438_store_0_req_1); -- 
    cr_1596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => type_cast_446_inst_req_1); -- 
    cr_2066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_load_1_req_1); -- 
    cr_2071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_load_2_req_1); -- 
    cr_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => ptr_deref_513_load_3_req_1); -- 
    cr_2095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(284), ack => type_cast_527_inst_req_1); -- 
    -- CP-element group 285:  transition  output  delay-element  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	212 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	289 
    -- CP-element group 285:  members (5) 
      -- CP-element group 285: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27_PhiReq/$exit
      -- CP-element group 285: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27_PhiReq/phi_stmt_583/$exit
      -- CP-element group 285: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/$exit
      -- CP-element group 285: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_587_konst_delay_trans
      -- CP-element group 285: 	 branch_block_stmt_275/bbx_xnph_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_req
      -- 
    phi_stmt_583_req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_583_req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(285), ack => phi_stmt_583_req_0); -- 
    -- Element group testConfigure_CP_684_elements(285) is a control-delay.
    cp_element_285_delay: control_delay_element  generic map(name => " 285_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(212), ack => testConfigure_CP_684_elements(285), clk => clk, reset =>reset);
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	254 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/Sample/ra
      -- 
    ra_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_589_inst_ack_0, ack => testConfigure_CP_684_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	254 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (2) 
      -- CP-element group 287: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/Update/ca
      -- 
    ca_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_589_inst_ack_1, ack => testConfigure_CP_684_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/$exit
      -- CP-element group 288: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/$exit
      -- CP-element group 288: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/$exit
      -- CP-element group 288: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/$exit
      -- CP-element group 288: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_589/SplitProtocol/$exit
      -- CP-element group 288: 	 branch_block_stmt_275/forx_xbody27_forx_xbody27_PhiReq/phi_stmt_583/phi_stmt_583_req
      -- 
    phi_stmt_583_req_2735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_583_req_2735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(288), ack => phi_stmt_583_req_1); -- 
    testConfigure_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(286) & testConfigure_CP_684_elements(287);
      gj_testConfigure_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  merge  transition  place  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	285 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (2) 
      -- CP-element group 289: 	 branch_block_stmt_275/merge_stmt_582_PhiReqMerge
      -- CP-element group 289: 	 branch_block_stmt_275/merge_stmt_582_PhiAck/$entry
      -- 
    testConfigure_CP_684_elements(289) <= OrReduce(testConfigure_CP_684_elements(285) & testConfigure_CP_684_elements(288));
    -- CP-element group 290:  fork  transition  place  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	213 
    -- CP-element group 290: 	214 
    -- CP-element group 290: 	216 
    -- CP-element group 290: 	217 
    -- CP-element group 290: 	220 
    -- CP-element group 290: 	224 
    -- CP-element group 290: 	228 
    -- CP-element group 290: 	232 
    -- CP-element group 290: 	236 
    -- CP-element group 290: 	240 
    -- CP-element group 290: 	244 
    -- CP-element group 290: 	248 
    -- CP-element group 290: 	251 
    -- CP-element group 290:  members (56) 
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745__entry__
      -- CP-element group 290: 	 branch_block_stmt_275/merge_stmt_582__exit__
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_resized_1
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_scaled_1
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_computed_1
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_resize_1/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_resize_1/$exit
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_resize_1/index_resize_req
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_resize_1/index_resize_ack
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_scale_1/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_scale_1/$exit
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_scale_1/scale_rename_req
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_index_scale_1/scale_rename_ack
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_update_start
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/array_obj_ref_595_final_index_sum_regn_Update/req
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_complete/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/addr_of_596_complete/req
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/RPIPE_zeropad_input_pipe_599_Sample/rr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_603_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_616_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_634_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_652_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_670_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_688_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_706_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/type_cast_724_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_update_start_
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Update/word_access_complete/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Update/word_access_complete/word_0/$entry
      -- CP-element group 290: 	 branch_block_stmt_275/assign_stmt_597_to_assign_stmt_745/ptr_deref_732_Update/word_access_complete/word_0/cr
      -- CP-element group 290: 	 branch_block_stmt_275/merge_stmt_582_PhiAck/$exit
      -- CP-element group 290: 	 branch_block_stmt_275/merge_stmt_582_PhiAck/phi_stmt_583_ack
      -- 
    phi_stmt_583_ack_2740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_583_ack_0, ack => testConfigure_CP_684_elements(290)); -- 
    req_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => array_obj_ref_595_index_offset_req_0); -- 
    req_2167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => array_obj_ref_595_index_offset_req_1); -- 
    req_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => addr_of_596_final_reg_req_1); -- 
    rr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => RPIPE_zeropad_input_pipe_599_inst_req_0); -- 
    cr_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => type_cast_603_inst_req_1); -- 
    cr_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => type_cast_616_inst_req_1); -- 
    cr_2266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => type_cast_634_inst_req_1); -- 
    cr_2294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => type_cast_652_inst_req_1); -- 
    cr_2322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => type_cast_670_inst_req_1); -- 
    cr_2350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => type_cast_688_inst_req_1); -- 
    cr_2378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => type_cast_706_inst_req_1); -- 
    cr_2406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => type_cast_724_inst_req_1); -- 
    cr_2456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(290), ack => ptr_deref_732_store_0_req_1); -- 
    -- CP-element group 291:  merge  fork  transition  place  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	209 
    -- CP-element group 291: 	253 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	255 
    -- CP-element group 291: 	256 
    -- CP-element group 291:  members (13) 
      -- CP-element group 291: 	 branch_block_stmt_275/merge_stmt_754_PhiAck/$exit
      -- CP-element group 291: 	 branch_block_stmt_275/merge_stmt_754_PhiAck/dummy
      -- CP-element group 291: 	 branch_block_stmt_275/assign_stmt_758__entry__
      -- CP-element group 291: 	 branch_block_stmt_275/merge_stmt_754__exit__
      -- CP-element group 291: 	 branch_block_stmt_275/merge_stmt_754_PhiAck/$entry
      -- CP-element group 291: 	 branch_block_stmt_275/assign_stmt_758/$entry
      -- CP-element group 291: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_sample_start_
      -- CP-element group 291: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_update_start_
      -- CP-element group 291: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_Sample/$entry
      -- CP-element group 291: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_Sample/rr
      -- CP-element group 291: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_275/assign_stmt_758/type_cast_757_Update/cr
      -- CP-element group 291: 	 branch_block_stmt_275/merge_stmt_754_PhiReqMerge
      -- 
    rr_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(291), ack => type_cast_757_inst_req_0); -- 
    cr_2492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(291), ack => type_cast_757_inst_req_1); -- 
    testConfigure_CP_684_elements(291) <= OrReduce(testConfigure_CP_684_elements(209) & testConfigure_CP_684_elements(253));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar96_362_resized : std_logic_vector(8 downto 0);
    signal R_indvar96_362_scaled : std_logic_vector(8 downto 0);
    signal R_indvar_594_resized : std_logic_vector(13 downto 0);
    signal R_indvar_594_scaled : std_logic_vector(13 downto 0);
    signal STORE_pad_419_data_0 : std_logic_vector(7 downto 0);
    signal STORE_pad_419_word_address_0 : std_logic_vector(0 downto 0);
    signal add40_640 : std_logic_vector(63 downto 0);
    signal add46_658 : std_logic_vector(63 downto 0);
    signal add52_676 : std_logic_vector(63 downto 0);
    signal add58_694 : std_logic_vector(63 downto 0);
    signal add64_712 : std_logic_vector(63 downto 0);
    signal add70_730 : std_logic_vector(63 downto 0);
    signal add_622 : std_logic_vector(63 downto 0);
    signal array_obj_ref_363_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_363_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_363_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_363_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_363_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_363_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_595_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_595_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_595_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_595_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_595_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_595_root_address : std_logic_vector(13 downto 0);
    signal arrayidx74_597 : std_logic_vector(31 downto 0);
    signal arrayidx_365 : std_logic_vector(31 downto 0);
    signal call11_443 : std_logic_vector(7 downto 0);
    signal call13_462 : std_logic_vector(7 downto 0);
    signal call1_302 : std_logic_vector(7 downto 0);
    signal call29_600 : std_logic_vector(7 downto 0);
    signal call32_613 : std_logic_vector(7 downto 0);
    signal call37_631 : std_logic_vector(7 downto 0);
    signal call43_649 : std_logic_vector(7 downto 0);
    signal call487_325 : std_logic_vector(7 downto 0);
    signal call489_342 : std_logic_vector(7 downto 0);
    signal call49_667 : std_logic_vector(7 downto 0);
    signal call4_397 : std_logic_vector(7 downto 0);
    signal call4x_xlcssa1_405 : std_logic_vector(7 downto 0);
    signal call4x_xlcssa_412 : std_logic_vector(7 downto 0);
    signal call55_685 : std_logic_vector(7 downto 0);
    signal call61_703 : std_logic_vector(7 downto 0);
    signal call67_721 : std_logic_vector(7 downto 0);
    signal call9_424 : std_logic_vector(7 downto 0);
    signal call_289 : std_logic_vector(7 downto 0);
    signal cmp2583_540 : std_logic_vector(0 downto 0);
    signal cmp86_322 : std_logic_vector(0 downto 0);
    signal cmp_394 : std_logic_vector(0 downto 0);
    signal conv10_428 : std_logic_vector(31 downto 0);
    signal conv12_447 : std_logic_vector(31 downto 0);
    signal conv14_466 : std_logic_vector(31 downto 0);
    signal conv20_528 : std_logic_vector(63 downto 0);
    signal conv30_604 : std_logic_vector(63 downto 0);
    signal conv34_617 : std_logic_vector(63 downto 0);
    signal conv39_635 : std_logic_vector(63 downto 0);
    signal conv45_653 : std_logic_vector(63 downto 0);
    signal conv51_671 : std_logic_vector(63 downto 0);
    signal conv57_689 : std_logic_vector(63 downto 0);
    signal conv5_369 : std_logic_vector(31 downto 0);
    signal conv63_707 : std_logic_vector(63 downto 0);
    signal conv69_725 : std_logic_vector(63 downto 0);
    signal conv_306 : std_logic_vector(31 downto 0);
    signal exitcond10_745 : std_logic_vector(0 downto 0);
    signal iNsTr_0_281 : std_logic_vector(31 downto 0);
    signal iNsTr_12_436 : std_logic_vector(31 downto 0);
    signal iNsTr_15_455 : std_logic_vector(31 downto 0);
    signal iNsTr_18_474 : std_logic_vector(31 downto 0);
    signal iNsTr_20_486 : std_logic_vector(31 downto 0);
    signal iNsTr_21_498 : std_logic_vector(31 downto 0);
    signal iNsTr_22_510 : std_logic_vector(31 downto 0);
    signal iNsTr_28_385 : std_logic_vector(31 downto 0);
    signal iNsTr_3_295 : std_logic_vector(31 downto 0);
    signal iNsTr_6_312 : std_logic_vector(31 downto 0);
    signal inc_358 : std_logic_vector(31 downto 0);
    signal indvar96_335 : std_logic_vector(63 downto 0);
    signal indvar_583 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_740 : std_logic_vector(63 downto 0);
    signal mul19_524 : std_logic_vector(31 downto 0);
    signal mul_519 : std_logic_vector(31 downto 0);
    signal ptr_deref_283_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_283_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_283_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_283_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_283_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_283_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_283_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_283_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_283_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_283_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_283_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_283_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_283_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_283_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_283_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_297_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_297_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_297_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_297_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_297_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_297_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_314_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_314_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_314_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_314_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_314_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_314_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_314_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_314_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_314_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_314_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_314_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_314_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_314_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_314_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_314_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_371_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_371_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_371_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_371_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_371_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_371_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_371_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_371_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_371_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_371_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_371_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_371_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_371_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_371_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_371_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_388_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_388_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_388_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_388_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_388_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_388_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_388_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_388_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_388_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_388_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_388_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_388_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_388_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_388_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_438_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_438_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_438_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_438_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_438_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_438_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_457_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_457_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_457_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_457_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_457_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_457_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_476_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_476_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_476_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_476_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_476_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_476_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_489_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_489_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_489_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_489_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_489_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_489_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_489_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_489_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_489_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_489_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_489_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_489_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_489_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_489_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_501_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_501_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_501_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_501_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_501_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_501_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_501_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_501_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_501_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_501_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_501_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_501_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_501_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_501_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_513_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_513_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_513_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_513_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_513_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_513_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_513_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_513_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_513_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_513_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_513_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_513_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_513_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_513_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_732_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_732_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_732_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_732_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_732_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_732_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl36_628 : std_logic_vector(63 downto 0);
    signal shl42_646 : std_logic_vector(63 downto 0);
    signal shl48_664 : std_logic_vector(63 downto 0);
    signal shl54_682 : std_logic_vector(63 downto 0);
    signal shl60_700 : std_logic_vector(63 downto 0);
    signal shl66_718 : std_logic_vector(63 downto 0);
    signal shl_610 : std_logic_vector(63 downto 0);
    signal shr82x_xmask_534 : std_logic_vector(63 downto 0);
    signal tmp16_490 : std_logic_vector(31 downto 0);
    signal tmp17_502 : std_logic_vector(31 downto 0);
    signal tmp18_514 : std_logic_vector(31 downto 0);
    signal tmp2_389 : std_logic_vector(31 downto 0);
    signal tmp4_552 : std_logic_vector(31 downto 0);
    signal tmp5_557 : std_logic_vector(31 downto 0);
    signal tmp6_561 : std_logic_vector(63 downto 0);
    signal tmp7_567 : std_logic_vector(63 downto 0);
    signal tmp8_573 : std_logic_vector(0 downto 0);
    signal tmp98_379 : std_logic_vector(63 downto 0);
    signal tmp_354 : std_logic_vector(63 downto 0);
    signal type_cast_285_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_320_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_338_wire : std_logic_vector(63 downto 0);
    signal type_cast_341_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_345_wire : std_logic_vector(7 downto 0);
    signal type_cast_347_wire : std_logic_vector(7 downto 0);
    signal type_cast_352_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_377_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_408_wire : std_logic_vector(7 downto 0);
    signal type_cast_415_wire : std_logic_vector(7 downto 0);
    signal type_cast_417_wire : std_logic_vector(7 downto 0);
    signal type_cast_532_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_538_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_565_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_571_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_578_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_587_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_589_wire : std_logic_vector(63 downto 0);
    signal type_cast_608_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_644_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_662_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_680_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_698_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_716_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(63 downto 0);
    signal umax9_580 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_pad_419_word_address_0 <= "0";
    array_obj_ref_363_constant_part_of_offset <= "000001001";
    array_obj_ref_363_offset_scale_factor_0 <= "100000000";
    array_obj_ref_363_offset_scale_factor_1 <= "000000100";
    array_obj_ref_363_resized_base_address <= "000000000";
    array_obj_ref_595_constant_part_of_offset <= "00000000000000";
    array_obj_ref_595_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_595_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_595_resized_base_address <= "00000000000000";
    iNsTr_0_281 <= "00000000000000000000000000000000";
    iNsTr_12_436 <= "00000000000000000000000000000010";
    iNsTr_15_455 <= "00000000000000000000000000000011";
    iNsTr_18_474 <= "00000000000000000000000000000100";
    iNsTr_20_486 <= "00000000000000000000000000001001";
    iNsTr_21_498 <= "00000000000000000000000000001101";
    iNsTr_22_510 <= "00000000000000000000000000010001";
    iNsTr_28_385 <= "00000000000000000000000000000101";
    iNsTr_3_295 <= "00000000000000000000000000000100";
    iNsTr_6_312 <= "00000000000000000000000000000101";
    ptr_deref_283_word_offset_0 <= "000000000";
    ptr_deref_283_word_offset_1 <= "000000001";
    ptr_deref_283_word_offset_2 <= "000000010";
    ptr_deref_283_word_offset_3 <= "000000011";
    ptr_deref_297_word_offset_0 <= "000000000";
    ptr_deref_314_word_offset_0 <= "000000000";
    ptr_deref_314_word_offset_1 <= "000000001";
    ptr_deref_314_word_offset_2 <= "000000010";
    ptr_deref_314_word_offset_3 <= "000000011";
    ptr_deref_371_word_offset_0 <= "000000000";
    ptr_deref_371_word_offset_1 <= "000000001";
    ptr_deref_371_word_offset_2 <= "000000010";
    ptr_deref_371_word_offset_3 <= "000000011";
    ptr_deref_388_word_offset_0 <= "000000000";
    ptr_deref_388_word_offset_1 <= "000000001";
    ptr_deref_388_word_offset_2 <= "000000010";
    ptr_deref_388_word_offset_3 <= "000000011";
    ptr_deref_438_word_offset_0 <= "0000000";
    ptr_deref_457_word_offset_0 <= "0000000";
    ptr_deref_476_word_offset_0 <= "0000000";
    ptr_deref_489_word_offset_0 <= "000000000";
    ptr_deref_489_word_offset_1 <= "000000001";
    ptr_deref_489_word_offset_2 <= "000000010";
    ptr_deref_489_word_offset_3 <= "000000011";
    ptr_deref_501_word_offset_0 <= "000000000";
    ptr_deref_501_word_offset_1 <= "000000001";
    ptr_deref_501_word_offset_2 <= "000000010";
    ptr_deref_501_word_offset_3 <= "000000011";
    ptr_deref_513_word_offset_0 <= "000000000";
    ptr_deref_513_word_offset_1 <= "000000001";
    ptr_deref_513_word_offset_2 <= "000000010";
    ptr_deref_513_word_offset_3 <= "000000011";
    ptr_deref_732_word_offset_0 <= "00000000000000";
    type_cast_285_wire_constant <= "00000000000000000000000000000101";
    type_cast_320_wire_constant <= "00000000";
    type_cast_341_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_352_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_377_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_532_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_538_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_565_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_571_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_578_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_587_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_608_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_626_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_644_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_662_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_680_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_698_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_716_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_738_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_335: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_338_wire & type_cast_341_wire_constant;
      req <= phi_stmt_335_req_0 & phi_stmt_335_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_335",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_335_ack_0,
          idata => idata,
          odata => indvar96_335,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_335
    phi_stmt_342: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_345_wire & type_cast_347_wire;
      req <= phi_stmt_342_req_0 & phi_stmt_342_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_342",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_342_ack_0,
          idata => idata,
          odata => call489_342,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_342
    phi_stmt_405: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_408_wire;
      req(0) <= phi_stmt_405_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_405",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_405_ack_0,
          idata => idata,
          odata => call4x_xlcssa1_405,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_405
    phi_stmt_412: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_415_wire & type_cast_417_wire;
      req <= phi_stmt_412_req_0 & phi_stmt_412_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_412",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_412_ack_0,
          idata => idata,
          odata => call4x_xlcssa_412,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_412
    phi_stmt_583: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_587_wire_constant & type_cast_589_wire;
      req <= phi_stmt_583_req_0 & phi_stmt_583_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_583",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_583_ack_0,
          idata => idata,
          odata => indvar_583,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_583
    -- flow-through select operator MUX_579_inst
    umax9_580 <= tmp7_567 when (tmp8_573(0) /=  '0') else type_cast_578_wire_constant;
    addr_of_364_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_364_final_reg_req_0;
      addr_of_364_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_364_final_reg_req_1;
      addr_of_364_final_reg_ack_1<= rack(0);
      addr_of_364_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_364_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 9,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_363_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_596_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_596_final_reg_req_0;
      addr_of_596_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_596_final_reg_req_1;
      addr_of_596_final_reg_ack_1<= rack(0);
      addr_of_596_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_596_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_595_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx74_597,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_305_inst_req_0;
      type_cast_305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_305_inst_req_1;
      type_cast_305_inst_ack_1<= rack(0);
      type_cast_305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_302,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_338_inst_req_0;
      type_cast_338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_338_inst_req_1;
      type_cast_338_inst_ack_1<= rack(0);
      type_cast_338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp98_379,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_338_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_345_inst_req_0;
      type_cast_345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_345_inst_req_1;
      type_cast_345_inst_ack_1<= rack(0);
      type_cast_345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_397,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_345_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_347_inst_req_0;
      type_cast_347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_347_inst_req_1;
      type_cast_347_inst_ack_1<= rack(0);
      type_cast_347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call487_325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_347_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_357_inst_req_0;
      type_cast_357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_357_inst_req_1;
      type_cast_357_inst_ack_1<= rack(0);
      type_cast_357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_368_inst_req_0;
      type_cast_368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_368_inst_req_1;
      type_cast_368_inst_ack_1<= rack(0);
      type_cast_368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call489_342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5_369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_408_inst_req_0;
      type_cast_408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_408_inst_req_1;
      type_cast_408_inst_ack_1<= rack(0);
      type_cast_408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_397,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_408_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_415_inst_req_0;
      type_cast_415_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_415_inst_req_1;
      type_cast_415_inst_ack_1<= rack(0);
      type_cast_415_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_415_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call487_325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_415_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_417_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_417_inst_req_0;
      type_cast_417_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_417_inst_req_1;
      type_cast_417_inst_ack_1<= rack(0);
      type_cast_417_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_417_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4x_xlcssa1_405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_417_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_427_inst_req_0;
      type_cast_427_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_427_inst_req_1;
      type_cast_427_inst_ack_1<= rack(0);
      type_cast_427_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_427_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call9_424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_446_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_446_inst_req_0;
      type_cast_446_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_446_inst_req_1;
      type_cast_446_inst_ack_1<= rack(0);
      type_cast_446_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_446_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_443,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_447,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_465_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_465_inst_req_0;
      type_cast_465_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_465_inst_req_1;
      type_cast_465_inst_ack_1<= rack(0);
      type_cast_465_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_465_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call13_462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_466,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_527_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_527_inst_req_0;
      type_cast_527_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_527_inst_req_1;
      type_cast_527_inst_ack_1<= rack(0);
      type_cast_527_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_527_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul19_524,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_528,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_560_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_560_inst_req_0;
      type_cast_560_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_560_inst_req_1;
      type_cast_560_inst_ack_1<= rack(0);
      type_cast_560_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_560_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_557,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_561,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_589_inst_req_0;
      type_cast_589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_589_inst_req_1;
      type_cast_589_inst_ack_1<= rack(0);
      type_cast_589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_740,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_589_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_603_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_603_inst_req_0;
      type_cast_603_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_603_inst_req_1;
      type_cast_603_inst_ack_1<= rack(0);
      type_cast_603_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_603_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29_600,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_604,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_616_inst_req_0;
      type_cast_616_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_616_inst_req_1;
      type_cast_616_inst_ack_1<= rack(0);
      type_cast_616_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_616_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_617,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_634_inst_req_0;
      type_cast_634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_634_inst_req_1;
      type_cast_634_inst_ack_1<= rack(0);
      type_cast_634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_652_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_652_inst_req_0;
      type_cast_652_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_652_inst_req_1;
      type_cast_652_inst_ack_1<= rack(0);
      type_cast_652_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_652_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call43_649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_653,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_670_inst_req_0;
      type_cast_670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_670_inst_req_1;
      type_cast_670_inst_ack_1<= rack(0);
      type_cast_670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call49_667,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_688_inst_req_0;
      type_cast_688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_688_inst_req_1;
      type_cast_688_inst_ack_1<= rack(0);
      type_cast_688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_685,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv57_689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_706_inst_req_0;
      type_cast_706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_706_inst_req_1;
      type_cast_706_inst_ack_1<= rack(0);
      type_cast_706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_707,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_724_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_724_inst_req_0;
      type_cast_724_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_724_inst_req_1;
      type_cast_724_inst_ack_1<= rack(0);
      type_cast_724_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_724_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call67_721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_725,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_757_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_757_inst_req_0;
      type_cast_757_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_757_inst_req_1;
      type_cast_757_inst_ack_1<= rack(0);
      type_cast_757_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_757_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul19_524,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_pad_419_gather_scatter
    process(call4x_xlcssa_412) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call4x_xlcssa_412;
      ov(7 downto 0) := iv;
      STORE_pad_419_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_363_index_1_resize
    process(indvar96_335) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar96_335;
      ov := iv(8 downto 0);
      R_indvar96_362_resized <= ov(8 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_363_root_address_inst
    process(array_obj_ref_363_final_offset) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_363_final_offset;
      ov(8 downto 0) := iv;
      array_obj_ref_363_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_595_index_1_rename
    process(R_indvar_594_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_594_resized;
      ov(13 downto 0) := iv;
      R_indvar_594_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_595_index_1_resize
    process(indvar_583) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_583;
      ov := iv(13 downto 0);
      R_indvar_594_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_595_root_address_inst
    process(array_obj_ref_595_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_595_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_595_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_283_base_resize
    process(iNsTr_0_281) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_281;
      ov := iv(8 downto 0);
      ptr_deref_283_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_283_gather_scatter
    process(type_cast_285_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_285_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_283_data_3 <= ov(31 downto 24);
      ptr_deref_283_data_2 <= ov(23 downto 16);
      ptr_deref_283_data_1 <= ov(15 downto 8);
      ptr_deref_283_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_283_root_address_inst
    process(ptr_deref_283_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_283_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_283_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_297_addr_0
    process(ptr_deref_297_root_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_297_root_address;
      ov(8 downto 0) := iv;
      ptr_deref_297_word_address_0 <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_297_base_resize
    process(iNsTr_3_295) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_295;
      ov := iv(8 downto 0);
      ptr_deref_297_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_297_gather_scatter
    process(call_289) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call_289;
      ov(7 downto 0) := iv;
      ptr_deref_297_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_297_root_address_inst
    process(ptr_deref_297_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_297_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_297_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_314_base_resize
    process(iNsTr_6_312) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_312;
      ov := iv(8 downto 0);
      ptr_deref_314_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_314_gather_scatter
    process(conv_306) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_306;
      ov(31 downto 0) := iv;
      ptr_deref_314_data_3 <= ov(31 downto 24);
      ptr_deref_314_data_2 <= ov(23 downto 16);
      ptr_deref_314_data_1 <= ov(15 downto 8);
      ptr_deref_314_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_314_root_address_inst
    process(ptr_deref_314_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_314_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_314_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_371_base_resize
    process(arrayidx_365) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_365;
      ov := iv(8 downto 0);
      ptr_deref_371_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_371_gather_scatter
    process(conv5_369) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv5_369;
      ov(31 downto 0) := iv;
      ptr_deref_371_data_3 <= ov(31 downto 24);
      ptr_deref_371_data_2 <= ov(23 downto 16);
      ptr_deref_371_data_1 <= ov(15 downto 8);
      ptr_deref_371_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_371_root_address_inst
    process(ptr_deref_371_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_371_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_371_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_388_base_resize
    process(iNsTr_28_385) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_28_385;
      ov := iv(8 downto 0);
      ptr_deref_388_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_388_gather_scatter
    process(ptr_deref_388_data_3, ptr_deref_388_data_2, ptr_deref_388_data_1, ptr_deref_388_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_388_data_3 & ptr_deref_388_data_2 & ptr_deref_388_data_1 & ptr_deref_388_data_0;
      ov(31 downto 0) := iv;
      tmp2_389 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_388_root_address_inst
    process(ptr_deref_388_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_388_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_388_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_addr_0
    process(ptr_deref_438_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_438_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_438_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_base_resize
    process(iNsTr_12_436) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_12_436;
      ov := iv(6 downto 0);
      ptr_deref_438_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_gather_scatter
    process(conv10_428) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv10_428;
      ov(31 downto 0) := iv;
      ptr_deref_438_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_root_address_inst
    process(ptr_deref_438_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_438_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_438_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_457_addr_0
    process(ptr_deref_457_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_457_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_457_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_457_base_resize
    process(iNsTr_15_455) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_15_455;
      ov := iv(6 downto 0);
      ptr_deref_457_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_457_gather_scatter
    process(conv12_447) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv12_447;
      ov(31 downto 0) := iv;
      ptr_deref_457_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_457_root_address_inst
    process(ptr_deref_457_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_457_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_457_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_476_addr_0
    process(ptr_deref_476_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_476_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_476_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_476_base_resize
    process(iNsTr_18_474) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_18_474;
      ov := iv(6 downto 0);
      ptr_deref_476_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_476_gather_scatter
    process(conv14_466) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv14_466;
      ov(31 downto 0) := iv;
      ptr_deref_476_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_476_root_address_inst
    process(ptr_deref_476_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_476_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_476_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_489_base_resize
    process(iNsTr_20_486) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_20_486;
      ov := iv(8 downto 0);
      ptr_deref_489_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_489_gather_scatter
    process(ptr_deref_489_data_3, ptr_deref_489_data_2, ptr_deref_489_data_1, ptr_deref_489_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_489_data_3 & ptr_deref_489_data_2 & ptr_deref_489_data_1 & ptr_deref_489_data_0;
      ov(31 downto 0) := iv;
      tmp16_490 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_489_root_address_inst
    process(ptr_deref_489_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_489_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_489_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_501_base_resize
    process(iNsTr_21_498) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_498;
      ov := iv(8 downto 0);
      ptr_deref_501_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_501_gather_scatter
    process(ptr_deref_501_data_3, ptr_deref_501_data_2, ptr_deref_501_data_1, ptr_deref_501_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_501_data_3 & ptr_deref_501_data_2 & ptr_deref_501_data_1 & ptr_deref_501_data_0;
      ov(31 downto 0) := iv;
      tmp17_502 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_501_root_address_inst
    process(ptr_deref_501_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_501_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_501_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_513_base_resize
    process(iNsTr_22_510) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_22_510;
      ov := iv(8 downto 0);
      ptr_deref_513_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_513_gather_scatter
    process(ptr_deref_513_data_3, ptr_deref_513_data_2, ptr_deref_513_data_1, ptr_deref_513_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_513_data_3 & ptr_deref_513_data_2 & ptr_deref_513_data_1 & ptr_deref_513_data_0;
      ov(31 downto 0) := iv;
      tmp18_514 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_513_root_address_inst
    process(ptr_deref_513_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_513_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_513_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_732_addr_0
    process(ptr_deref_732_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_732_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_732_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_732_base_resize
    process(arrayidx74_597) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx74_597;
      ov := iv(13 downto 0);
      ptr_deref_732_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_732_gather_scatter
    process(add70_730) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add70_730;
      ov(63 downto 0) := iv;
      ptr_deref_732_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_732_root_address_inst
    process(ptr_deref_732_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_732_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_732_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_326_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp86_322;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_326_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_326_branch_req_0,
          ack0 => if_stmt_326_branch_ack_0,
          ack1 => if_stmt_326_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_398_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_394;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_398_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_398_branch_req_0,
          ack0 => if_stmt_398_branch_ack_0,
          ack1 => if_stmt_398_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_541_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp2583_540;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_541_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_541_branch_req_0,
          ack0 => if_stmt_541_branch_ack_0,
          ack1 => if_stmt_541_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_746_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond10_745;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_746_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_746_branch_req_0,
          ack0 => if_stmt_746_branch_ack_0,
          ack1 => if_stmt_746_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_353_inst
    process(indvar96_335) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar96_335, type_cast_352_wire_constant, tmp_var);
      tmp_354 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_378_inst
    process(indvar96_335) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar96_335, type_cast_377_wire_constant, tmp_var);
      tmp98_379 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_739_inst
    process(indvar_583) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_583, type_cast_738_wire_constant, tmp_var);
      indvarx_xnext_740 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_533_inst
    process(conv20_528) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv20_528, type_cast_532_wire_constant, tmp_var);
      shr82x_xmask_534 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_539_inst
    process(shr82x_xmask_534) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr82x_xmask_534, type_cast_538_wire_constant, tmp_var);
      cmp2583_540 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_744_inst
    process(indvarx_xnext_740, umax9_580) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_740, umax9_580, tmp_var);
      exitcond10_745 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_321_inst
    process(call1_302) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(call1_302, type_cast_320_wire_constant, tmp_var);
      cmp86_322 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_566_inst
    process(tmp6_561) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp6_561, type_cast_565_wire_constant, tmp_var);
      tmp7_567 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_518_inst
    process(tmp17_502, tmp16_490) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp17_502, tmp16_490, tmp_var);
      mul_519 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_523_inst
    process(mul_519, tmp18_514) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_519, tmp18_514, tmp_var);
      mul19_524 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_551_inst
    process(tmp17_502, tmp16_490) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp17_502, tmp16_490, tmp_var);
      tmp4_552 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_556_inst
    process(tmp4_552, tmp18_514) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp4_552, tmp18_514, tmp_var);
      tmp5_557 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_621_inst
    process(shl_610, conv34_617) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_610, conv34_617, tmp_var);
      add_622 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_639_inst
    process(shl36_628, conv39_635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_628, conv39_635, tmp_var);
      add40_640 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_657_inst
    process(shl42_646, conv45_653) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl42_646, conv45_653, tmp_var);
      add46_658 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_675_inst
    process(shl48_664, conv51_671) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl48_664, conv51_671, tmp_var);
      add52_676 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_693_inst
    process(shl54_682, conv57_689) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_682, conv57_689, tmp_var);
      add58_694 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_711_inst
    process(shl60_700, conv63_707) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_700, conv63_707, tmp_var);
      add64_712 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_729_inst
    process(shl66_718, conv69_725) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl66_718, conv69_725, tmp_var);
      add70_730 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_609_inst
    process(conv30_604) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv30_604, type_cast_608_wire_constant, tmp_var);
      shl_610 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_627_inst
    process(add_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_622, type_cast_626_wire_constant, tmp_var);
      shl36_628 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_645_inst
    process(add40_640) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add40_640, type_cast_644_wire_constant, tmp_var);
      shl42_646 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_663_inst
    process(add46_658) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add46_658, type_cast_662_wire_constant, tmp_var);
      shl48_664 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_681_inst
    process(add52_676) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add52_676, type_cast_680_wire_constant, tmp_var);
      shl54_682 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_699_inst
    process(add58_694) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add58_694, type_cast_698_wire_constant, tmp_var);
      shl60_700 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_717_inst
    process(add64_712) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add64_712, type_cast_716_wire_constant, tmp_var);
      shl66_718 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_572_inst
    process(tmp7_567) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp7_567, type_cast_571_wire_constant, tmp_var);
      tmp8_573 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_393_inst
    process(inc_358, tmp2_389) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc_358, tmp2_389, tmp_var);
      cmp_394 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_363_index_1_scale 
    ApIntMul_group_28: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar96_362_resized;
      R_indvar96_362_scaled <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_363_index_1_scale_req_0;
      array_obj_ref_363_index_1_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_363_index_1_scale_req_1;
      array_obj_ref_363_index_1_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_28_gI: SplitGuardInterface generic map(name => "ApIntMul_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000100",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_363_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar96_362_scaled;
      array_obj_ref_363_final_offset <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_363_index_offset_req_0;
      array_obj_ref_363_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_363_index_offset_req_1;
      array_obj_ref_363_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000001001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_595_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_594_scaled;
      array_obj_ref_595_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_595_index_offset_req_0;
      array_obj_ref_595_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_595_index_offset_req_1;
      array_obj_ref_595_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : ptr_deref_283_addr_0 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_283_root_address;
      ptr_deref_283_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_283_addr_0_req_0;
      ptr_deref_283_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_283_addr_0_req_1;
      ptr_deref_283_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : ptr_deref_283_addr_1 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_283_root_address;
      ptr_deref_283_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_283_addr_1_req_0;
      ptr_deref_283_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_283_addr_1_req_1;
      ptr_deref_283_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : ptr_deref_283_addr_2 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_283_root_address;
      ptr_deref_283_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_283_addr_2_req_0;
      ptr_deref_283_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_283_addr_2_req_1;
      ptr_deref_283_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : ptr_deref_283_addr_3 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_283_root_address;
      ptr_deref_283_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_283_addr_3_req_0;
      ptr_deref_283_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_283_addr_3_req_1;
      ptr_deref_283_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : ptr_deref_314_addr_0 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_314_root_address;
      ptr_deref_314_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_314_addr_0_req_0;
      ptr_deref_314_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_314_addr_0_req_1;
      ptr_deref_314_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : ptr_deref_314_addr_1 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_314_root_address;
      ptr_deref_314_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_314_addr_1_req_0;
      ptr_deref_314_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_314_addr_1_req_1;
      ptr_deref_314_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : ptr_deref_314_addr_2 
    ApIntAdd_group_37: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_314_root_address;
      ptr_deref_314_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_314_addr_2_req_0;
      ptr_deref_314_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_314_addr_2_req_1;
      ptr_deref_314_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_37_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : ptr_deref_314_addr_3 
    ApIntAdd_group_38: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_314_root_address;
      ptr_deref_314_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_314_addr_3_req_0;
      ptr_deref_314_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_314_addr_3_req_1;
      ptr_deref_314_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_38_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : ptr_deref_371_addr_0 
    ApIntAdd_group_39: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_371_root_address;
      ptr_deref_371_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_371_addr_0_req_0;
      ptr_deref_371_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_371_addr_0_req_1;
      ptr_deref_371_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_39_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_39_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : ptr_deref_371_addr_1 
    ApIntAdd_group_40: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_371_root_address;
      ptr_deref_371_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_371_addr_1_req_0;
      ptr_deref_371_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_371_addr_1_req_1;
      ptr_deref_371_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_40_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_40_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_40",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : ptr_deref_371_addr_2 
    ApIntAdd_group_41: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_371_root_address;
      ptr_deref_371_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_371_addr_2_req_0;
      ptr_deref_371_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_371_addr_2_req_1;
      ptr_deref_371_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_41_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_41_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : ptr_deref_371_addr_3 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_371_root_address;
      ptr_deref_371_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_371_addr_3_req_0;
      ptr_deref_371_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_371_addr_3_req_1;
      ptr_deref_371_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : ptr_deref_388_addr_0 
    ApIntAdd_group_43: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_388_root_address;
      ptr_deref_388_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_388_addr_0_req_0;
      ptr_deref_388_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_388_addr_0_req_1;
      ptr_deref_388_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_43_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_43_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_43",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : ptr_deref_388_addr_1 
    ApIntAdd_group_44: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_388_root_address;
      ptr_deref_388_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_388_addr_1_req_0;
      ptr_deref_388_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_388_addr_1_req_1;
      ptr_deref_388_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_44_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_44_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : ptr_deref_388_addr_2 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_388_root_address;
      ptr_deref_388_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_388_addr_2_req_0;
      ptr_deref_388_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_388_addr_2_req_1;
      ptr_deref_388_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : ptr_deref_388_addr_3 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_388_root_address;
      ptr_deref_388_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_388_addr_3_req_0;
      ptr_deref_388_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_388_addr_3_req_1;
      ptr_deref_388_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : ptr_deref_489_addr_0 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_489_addr_0_req_0;
      ptr_deref_489_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_489_addr_0_req_1;
      ptr_deref_489_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : ptr_deref_489_addr_1 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_489_addr_1_req_0;
      ptr_deref_489_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_489_addr_1_req_1;
      ptr_deref_489_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : ptr_deref_489_addr_2 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_489_addr_2_req_0;
      ptr_deref_489_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_489_addr_2_req_1;
      ptr_deref_489_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : ptr_deref_489_addr_3 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_489_addr_3_req_0;
      ptr_deref_489_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_489_addr_3_req_1;
      ptr_deref_489_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : ptr_deref_501_addr_0 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_501_root_address;
      ptr_deref_501_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_501_addr_0_req_0;
      ptr_deref_501_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_501_addr_0_req_1;
      ptr_deref_501_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : ptr_deref_501_addr_1 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_501_root_address;
      ptr_deref_501_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_501_addr_1_req_0;
      ptr_deref_501_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_501_addr_1_req_1;
      ptr_deref_501_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : ptr_deref_501_addr_2 
    ApIntAdd_group_53: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_501_root_address;
      ptr_deref_501_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_501_addr_2_req_0;
      ptr_deref_501_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_501_addr_2_req_1;
      ptr_deref_501_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_53_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_53_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : ptr_deref_501_addr_3 
    ApIntAdd_group_54: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_501_root_address;
      ptr_deref_501_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_501_addr_3_req_0;
      ptr_deref_501_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_501_addr_3_req_1;
      ptr_deref_501_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_54_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_54_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_54",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : ptr_deref_513_addr_0 
    ApIntAdd_group_55: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_513_root_address;
      ptr_deref_513_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_513_addr_0_req_0;
      ptr_deref_513_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_513_addr_0_req_1;
      ptr_deref_513_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_55_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_55_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_55",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : ptr_deref_513_addr_1 
    ApIntAdd_group_56: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_513_root_address;
      ptr_deref_513_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_513_addr_1_req_0;
      ptr_deref_513_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_513_addr_1_req_1;
      ptr_deref_513_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_56_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_56_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_56",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : ptr_deref_513_addr_2 
    ApIntAdd_group_57: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_513_root_address;
      ptr_deref_513_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_513_addr_2_req_0;
      ptr_deref_513_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_513_addr_2_req_1;
      ptr_deref_513_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_57_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_57_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_57",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : ptr_deref_513_addr_3 
    ApIntAdd_group_58: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_513_root_address;
      ptr_deref_513_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_513_addr_3_req_0;
      ptr_deref_513_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_513_addr_3_req_1;
      ptr_deref_513_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_58_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_58_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_58",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared load operator group (0) : ptr_deref_388_load_0 ptr_deref_388_load_1 ptr_deref_388_load_2 ptr_deref_388_load_3 ptr_deref_489_load_0 ptr_deref_489_load_1 ptr_deref_489_load_2 ptr_deref_489_load_3 ptr_deref_501_load_0 ptr_deref_501_load_1 ptr_deref_501_load_2 ptr_deref_501_load_3 ptr_deref_513_load_0 ptr_deref_513_load_1 ptr_deref_513_load_2 ptr_deref_513_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(143 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_388_load_0_req_0;
      reqL_unguarded(14) <= ptr_deref_388_load_1_req_0;
      reqL_unguarded(13) <= ptr_deref_388_load_2_req_0;
      reqL_unguarded(12) <= ptr_deref_388_load_3_req_0;
      reqL_unguarded(11) <= ptr_deref_489_load_0_req_0;
      reqL_unguarded(10) <= ptr_deref_489_load_1_req_0;
      reqL_unguarded(9) <= ptr_deref_489_load_2_req_0;
      reqL_unguarded(8) <= ptr_deref_489_load_3_req_0;
      reqL_unguarded(7) <= ptr_deref_501_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_501_load_1_req_0;
      reqL_unguarded(5) <= ptr_deref_501_load_2_req_0;
      reqL_unguarded(4) <= ptr_deref_501_load_3_req_0;
      reqL_unguarded(3) <= ptr_deref_513_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_513_load_1_req_0;
      reqL_unguarded(1) <= ptr_deref_513_load_2_req_0;
      reqL_unguarded(0) <= ptr_deref_513_load_3_req_0;
      ptr_deref_388_load_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_388_load_1_ack_0 <= ackL_unguarded(14);
      ptr_deref_388_load_2_ack_0 <= ackL_unguarded(13);
      ptr_deref_388_load_3_ack_0 <= ackL_unguarded(12);
      ptr_deref_489_load_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_489_load_1_ack_0 <= ackL_unguarded(10);
      ptr_deref_489_load_2_ack_0 <= ackL_unguarded(9);
      ptr_deref_489_load_3_ack_0 <= ackL_unguarded(8);
      ptr_deref_501_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_501_load_1_ack_0 <= ackL_unguarded(6);
      ptr_deref_501_load_2_ack_0 <= ackL_unguarded(5);
      ptr_deref_501_load_3_ack_0 <= ackL_unguarded(4);
      ptr_deref_513_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_513_load_1_ack_0 <= ackL_unguarded(2);
      ptr_deref_513_load_2_ack_0 <= ackL_unguarded(1);
      ptr_deref_513_load_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_388_load_0_req_1;
      reqR_unguarded(14) <= ptr_deref_388_load_1_req_1;
      reqR_unguarded(13) <= ptr_deref_388_load_2_req_1;
      reqR_unguarded(12) <= ptr_deref_388_load_3_req_1;
      reqR_unguarded(11) <= ptr_deref_489_load_0_req_1;
      reqR_unguarded(10) <= ptr_deref_489_load_1_req_1;
      reqR_unguarded(9) <= ptr_deref_489_load_2_req_1;
      reqR_unguarded(8) <= ptr_deref_489_load_3_req_1;
      reqR_unguarded(7) <= ptr_deref_501_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_501_load_1_req_1;
      reqR_unguarded(5) <= ptr_deref_501_load_2_req_1;
      reqR_unguarded(4) <= ptr_deref_501_load_3_req_1;
      reqR_unguarded(3) <= ptr_deref_513_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_513_load_1_req_1;
      reqR_unguarded(1) <= ptr_deref_513_load_2_req_1;
      reqR_unguarded(0) <= ptr_deref_513_load_3_req_1;
      ptr_deref_388_load_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_388_load_1_ack_1 <= ackR_unguarded(14);
      ptr_deref_388_load_2_ack_1 <= ackR_unguarded(13);
      ptr_deref_388_load_3_ack_1 <= ackR_unguarded(12);
      ptr_deref_489_load_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_489_load_1_ack_1 <= ackR_unguarded(10);
      ptr_deref_489_load_2_ack_1 <= ackR_unguarded(9);
      ptr_deref_489_load_3_ack_1 <= ackR_unguarded(8);
      ptr_deref_501_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_501_load_1_ack_1 <= ackR_unguarded(6);
      ptr_deref_501_load_2_ack_1 <= ackR_unguarded(5);
      ptr_deref_501_load_3_ack_1 <= ackR_unguarded(4);
      ptr_deref_513_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_513_load_1_ack_1 <= ackR_unguarded(2);
      ptr_deref_513_load_2_ack_1 <= ackR_unguarded(1);
      ptr_deref_513_load_3_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_388_word_address_0 & ptr_deref_388_word_address_1 & ptr_deref_388_word_address_2 & ptr_deref_388_word_address_3 & ptr_deref_489_word_address_0 & ptr_deref_489_word_address_1 & ptr_deref_489_word_address_2 & ptr_deref_489_word_address_3 & ptr_deref_501_word_address_0 & ptr_deref_501_word_address_1 & ptr_deref_501_word_address_2 & ptr_deref_501_word_address_3 & ptr_deref_513_word_address_0 & ptr_deref_513_word_address_1 & ptr_deref_513_word_address_2 & ptr_deref_513_word_address_3;
      ptr_deref_388_data_0 <= data_out(127 downto 120);
      ptr_deref_388_data_1 <= data_out(119 downto 112);
      ptr_deref_388_data_2 <= data_out(111 downto 104);
      ptr_deref_388_data_3 <= data_out(103 downto 96);
      ptr_deref_489_data_0 <= data_out(95 downto 88);
      ptr_deref_489_data_1 <= data_out(87 downto 80);
      ptr_deref_489_data_2 <= data_out(79 downto 72);
      ptr_deref_489_data_3 <= data_out(71 downto 64);
      ptr_deref_501_data_0 <= data_out(63 downto 56);
      ptr_deref_501_data_1 <= data_out(55 downto 48);
      ptr_deref_501_data_2 <= data_out(47 downto 40);
      ptr_deref_501_data_3 <= data_out(39 downto 32);
      ptr_deref_513_data_0 <= data_out(31 downto 24);
      ptr_deref_513_data_1 <= data_out(23 downto 16);
      ptr_deref_513_data_2 <= data_out(15 downto 8);
      ptr_deref_513_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 9,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(8 downto 0),
          mtag => memory_space_2_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 16,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_pad_419_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_pad_419_store_0_req_0;
      STORE_pad_419_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_pad_419_store_0_req_1;
      STORE_pad_419_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_pad_419_word_address_0;
      data_in <= STORE_pad_419_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_314_store_1 ptr_deref_283_store_3 ptr_deref_314_store_0 ptr_deref_283_store_2 ptr_deref_297_store_0 ptr_deref_283_store_1 ptr_deref_283_store_0 ptr_deref_314_store_2 ptr_deref_314_store_3 ptr_deref_371_store_0 ptr_deref_371_store_1 ptr_deref_371_store_2 ptr_deref_371_store_3 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(116 downto 0);
      signal data_in: std_logic_vector(103 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 12 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 12 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant inBUFs : IntegerArray(12 downto 0) := (12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(12 downto 0) := (12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      reqL_unguarded(12) <= ptr_deref_314_store_1_req_0;
      reqL_unguarded(11) <= ptr_deref_283_store_3_req_0;
      reqL_unguarded(10) <= ptr_deref_314_store_0_req_0;
      reqL_unguarded(9) <= ptr_deref_283_store_2_req_0;
      reqL_unguarded(8) <= ptr_deref_297_store_0_req_0;
      reqL_unguarded(7) <= ptr_deref_283_store_1_req_0;
      reqL_unguarded(6) <= ptr_deref_283_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_314_store_2_req_0;
      reqL_unguarded(4) <= ptr_deref_314_store_3_req_0;
      reqL_unguarded(3) <= ptr_deref_371_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_371_store_1_req_0;
      reqL_unguarded(1) <= ptr_deref_371_store_2_req_0;
      reqL_unguarded(0) <= ptr_deref_371_store_3_req_0;
      ptr_deref_314_store_1_ack_0 <= ackL_unguarded(12);
      ptr_deref_283_store_3_ack_0 <= ackL_unguarded(11);
      ptr_deref_314_store_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_283_store_2_ack_0 <= ackL_unguarded(9);
      ptr_deref_297_store_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_283_store_1_ack_0 <= ackL_unguarded(7);
      ptr_deref_283_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_314_store_2_ack_0 <= ackL_unguarded(5);
      ptr_deref_314_store_3_ack_0 <= ackL_unguarded(4);
      ptr_deref_371_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_371_store_1_ack_0 <= ackL_unguarded(2);
      ptr_deref_371_store_2_ack_0 <= ackL_unguarded(1);
      ptr_deref_371_store_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(12) <= ptr_deref_314_store_1_req_1;
      reqR_unguarded(11) <= ptr_deref_283_store_3_req_1;
      reqR_unguarded(10) <= ptr_deref_314_store_0_req_1;
      reqR_unguarded(9) <= ptr_deref_283_store_2_req_1;
      reqR_unguarded(8) <= ptr_deref_297_store_0_req_1;
      reqR_unguarded(7) <= ptr_deref_283_store_1_req_1;
      reqR_unguarded(6) <= ptr_deref_283_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_314_store_2_req_1;
      reqR_unguarded(4) <= ptr_deref_314_store_3_req_1;
      reqR_unguarded(3) <= ptr_deref_371_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_371_store_1_req_1;
      reqR_unguarded(1) <= ptr_deref_371_store_2_req_1;
      reqR_unguarded(0) <= ptr_deref_371_store_3_req_1;
      ptr_deref_314_store_1_ack_1 <= ackR_unguarded(12);
      ptr_deref_283_store_3_ack_1 <= ackR_unguarded(11);
      ptr_deref_314_store_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_283_store_2_ack_1 <= ackR_unguarded(9);
      ptr_deref_297_store_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_283_store_1_ack_1 <= ackR_unguarded(7);
      ptr_deref_283_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_314_store_2_ack_1 <= ackR_unguarded(5);
      ptr_deref_314_store_3_ack_1 <= ackR_unguarded(4);
      ptr_deref_371_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_371_store_1_ack_1 <= ackR_unguarded(2);
      ptr_deref_371_store_2_ack_1 <= ackR_unguarded(1);
      ptr_deref_371_store_3_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_11: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_12: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_314_word_address_1 & ptr_deref_283_word_address_3 & ptr_deref_314_word_address_0 & ptr_deref_283_word_address_2 & ptr_deref_297_word_address_0 & ptr_deref_283_word_address_1 & ptr_deref_283_word_address_0 & ptr_deref_314_word_address_2 & ptr_deref_314_word_address_3 & ptr_deref_371_word_address_0 & ptr_deref_371_word_address_1 & ptr_deref_371_word_address_2 & ptr_deref_371_word_address_3;
      data_in <= ptr_deref_314_data_1 & ptr_deref_283_data_3 & ptr_deref_314_data_0 & ptr_deref_283_data_2 & ptr_deref_297_data_0 & ptr_deref_283_data_1 & ptr_deref_283_data_0 & ptr_deref_314_data_2 & ptr_deref_314_data_3 & ptr_deref_371_data_0 & ptr_deref_371_data_1 & ptr_deref_371_data_2 & ptr_deref_371_data_3;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 9,
        data_width => 8,
        num_reqs => 13,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(8 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 13,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_438_store_0 ptr_deref_457_store_0 ptr_deref_476_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_438_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_457_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_476_store_0_req_0;
      ptr_deref_438_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_457_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_476_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_438_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_457_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_476_store_0_req_1;
      ptr_deref_438_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_457_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_476_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_438_word_address_0 & ptr_deref_457_word_address_0 & ptr_deref_476_word_address_0;
      data_in <= ptr_deref_438_data_0 & ptr_deref_457_data_0 & ptr_deref_476_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(6 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_732_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_732_store_0_req_0;
      ptr_deref_732_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_732_store_0_req_1;
      ptr_deref_732_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_732_word_address_0;
      data_in <= ptr_deref_732_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared inport operator group (0) : RPIPE_zeropad_input_pipe_301_inst RPIPE_zeropad_input_pipe_288_inst RPIPE_zeropad_input_pipe_324_inst RPIPE_zeropad_input_pipe_396_inst RPIPE_zeropad_input_pipe_423_inst RPIPE_zeropad_input_pipe_442_inst RPIPE_zeropad_input_pipe_461_inst RPIPE_zeropad_input_pipe_599_inst RPIPE_zeropad_input_pipe_612_inst RPIPE_zeropad_input_pipe_630_inst RPIPE_zeropad_input_pipe_648_inst RPIPE_zeropad_input_pipe_666_inst RPIPE_zeropad_input_pipe_684_inst RPIPE_zeropad_input_pipe_702_inst RPIPE_zeropad_input_pipe_720_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(119 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 14 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 14 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 14 downto 0);
      signal guard_vector : std_logic_vector( 14 downto 0);
      constant outBUFs : IntegerArray(14 downto 0) := (14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(14 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false);
      constant guardBuffering: IntegerArray(14 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2);
      -- 
    begin -- 
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_301_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_288_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_324_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_396_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_423_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_442_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_461_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_599_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_612_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_630_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_648_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_666_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_684_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_702_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_720_inst_req_0;
      RPIPE_zeropad_input_pipe_301_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_288_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_324_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_396_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_423_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_442_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_461_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_599_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_612_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_630_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_648_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_666_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_684_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_702_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_720_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_301_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_288_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_324_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_396_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_423_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_442_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_461_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_599_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_612_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_630_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_648_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_666_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_684_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_702_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_720_inst_req_1;
      RPIPE_zeropad_input_pipe_301_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_288_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_324_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_396_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_423_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_442_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_461_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_599_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_612_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_630_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_648_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_666_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_684_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_702_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_720_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      call1_302 <= data_out(119 downto 112);
      call_289 <= data_out(111 downto 104);
      call487_325 <= data_out(103 downto 96);
      call4_397 <= data_out(95 downto 88);
      call9_424 <= data_out(87 downto 80);
      call11_443 <= data_out(79 downto 72);
      call13_462 <= data_out(71 downto 64);
      call29_600 <= data_out(63 downto 56);
      call32_613 <= data_out(55 downto 48);
      call37_631 <= data_out(47 downto 40);
      call43_649 <= data_out(39 downto 32);
      call49_667 <= data_out(31 downto 24);
      call55_685 <= data_out(23 downto 16);
      call61_703 <= data_out(15 downto 8);
      call67_721 <= data_out(7 downto 0);
      zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_0_gI", nreqs => 15, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 15,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_2772_start: Boolean;
  signal zeropad3D_CP_2772_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_766_call_req_0 : boolean;
  signal call_stmt_766_call_ack_0 : boolean;
  signal call_stmt_766_call_req_1 : boolean;
  signal call_stmt_766_call_ack_1 : boolean;
  signal type_cast_770_inst_req_0 : boolean;
  signal type_cast_770_inst_ack_0 : boolean;
  signal type_cast_770_inst_req_1 : boolean;
  signal type_cast_770_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_772_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_772_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_772_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_772_inst_ack_1 : boolean;
  signal RPIPE_Block0_complete_776_inst_req_0 : boolean;
  signal RPIPE_Block0_complete_776_inst_ack_0 : boolean;
  signal RPIPE_Block0_complete_776_inst_req_1 : boolean;
  signal RPIPE_Block0_complete_776_inst_ack_1 : boolean;
  signal call_stmt_779_call_req_0 : boolean;
  signal call_stmt_779_call_ack_0 : boolean;
  signal call_stmt_779_call_req_1 : boolean;
  signal call_stmt_779_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_2772_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2772_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_2772_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2772_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_2772: Block -- control-path 
    signal zeropad3D_CP_2772_elements: BooleanArray(11 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_2772_elements(0) <= zeropad3D_CP_2772_start;
    zeropad3D_CP_2772_symbol <= zeropad3D_CP_2772_elements(11);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_764/$entry
      -- CP-element group 0: 	 branch_block_stmt_764/branch_block_stmt_764__entry__
      -- CP-element group 0: 	 branch_block_stmt_764/call_stmt_766__entry__
      -- CP-element group 0: 	 branch_block_stmt_764/call_stmt_766/$entry
      -- CP-element group 0: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_update_start_
      -- CP-element group 0: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_Update/ccr
      -- 
    crr_2798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(0), ack => call_stmt_766_call_req_0); -- 
    ccr_2803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(0), ack => call_stmt_766_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_Sample/cra
      -- 
    cra_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_766_call_ack_0, ack => zeropad3D_CP_2772_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (16) 
      -- CP-element group 2: 	 branch_block_stmt_764/call_stmt_766__exit__
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777__entry__
      -- CP-element group 2: 	 branch_block_stmt_764/call_stmt_766/$exit
      -- CP-element group 2: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_764/call_stmt_766/call_stmt_766_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/$entry
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_update_start_
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_Sample/rr
      -- 
    cca_2804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_766_call_ack_1, ack => zeropad3D_CP_2772_elements(2)); -- 
    rr_2815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(2), ack => type_cast_770_inst_req_0); -- 
    cr_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(2), ack => type_cast_770_inst_req_1); -- 
    rr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(2), ack => RPIPE_Block0_complete_776_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_Sample/ra
      -- 
    ra_2816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_770_inst_ack_0, ack => zeropad3D_CP_2772_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/type_cast_770_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_Sample/req
      -- 
    ca_2821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_770_inst_ack_1, ack => zeropad3D_CP_2772_elements(4)); -- 
    req_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(4), ack => WPIPE_Block0_starting_772_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_update_start_
      -- CP-element group 5: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_Update/req
      -- 
    ack_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_772_inst_ack_0, ack => zeropad3D_CP_2772_elements(5)); -- 
    req_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(5), ack => WPIPE_Block0_starting_772_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/WPIPE_Block0_starting_772_Update/ack
      -- 
    ack_2835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_772_inst_ack_1, ack => zeropad3D_CP_2772_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_update_start_
      -- CP-element group 7: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_Update/cr
      -- 
    ra_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_776_inst_ack_0, ack => zeropad3D_CP_2772_elements(7)); -- 
    cr_2848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(7), ack => RPIPE_Block0_complete_776_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/RPIPE_Block0_complete_776_Update/ca
      -- 
    ca_2849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_776_inst_ack_1, ack => zeropad3D_CP_2772_elements(8)); -- 
    -- CP-element group 9:  join  fork  transition  place  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777__exit__
      -- CP-element group 9: 	 branch_block_stmt_764/call_stmt_779__entry__
      -- CP-element group 9: 	 branch_block_stmt_764/assign_stmt_771_to_assign_stmt_777/$exit
      -- CP-element group 9: 	 branch_block_stmt_764/call_stmt_779/$entry
      -- CP-element group 9: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_update_start_
      -- CP-element group 9: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_Sample/crr
      -- CP-element group 9: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_Update/ccr
      -- 
    crr_2860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(9), ack => call_stmt_779_call_req_0); -- 
    ccr_2865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2772_elements(9), ack => call_stmt_779_call_req_1); -- 
    zeropad3D_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad3D_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2772_elements(6) & zeropad3D_CP_2772_elements(8);
      gj_zeropad3D_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2772_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_Sample/cra
      -- 
    cra_2861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_779_call_ack_0, ack => zeropad3D_CP_2772_elements(10)); -- 
    -- CP-element group 11:  transition  place  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (16) 
      -- CP-element group 11: 	 $exit
      -- CP-element group 11: 	 branch_block_stmt_764/$exit
      -- CP-element group 11: 	 branch_block_stmt_764/branch_block_stmt_764__exit__
      -- CP-element group 11: 	 branch_block_stmt_764/call_stmt_779__exit__
      -- CP-element group 11: 	 branch_block_stmt_764/return__
      -- CP-element group 11: 	 branch_block_stmt_764/merge_stmt_781__exit__
      -- CP-element group 11: 	 branch_block_stmt_764/call_stmt_779/$exit
      -- CP-element group 11: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_764/call_stmt_779/call_stmt_779_Update/cca
      -- CP-element group 11: 	 branch_block_stmt_764/return___PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_764/return___PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_764/merge_stmt_781_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_764/merge_stmt_781_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_764/merge_stmt_781_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_764/merge_stmt_781_PhiAck/dummy
      -- 
    cca_2866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_779_call_ack_1, ack => zeropad3D_CP_2772_elements(11)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call2_777 : std_logic_vector(7 downto 0);
    signal call_766 : std_logic_vector(15 downto 0);
    signal conv_771 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    type_cast_770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_770_inst_req_0;
      type_cast_770_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_770_inst_req_1;
      type_cast_770_inst_ack_1<= rack(0);
      type_cast_770_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_770_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_766,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_771,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- shared inport operator group (0) : RPIPE_Block0_complete_776_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_complete_776_inst_req_0;
      RPIPE_Block0_complete_776_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_complete_776_inst_req_1;
      RPIPE_Block0_complete_776_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call2_777 <= data_out(7 downto 0);
      Block0_complete_read_0_gI: SplitGuardInterface generic map(name => "Block0_complete_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_complete_read_0: InputPortRevised -- 
        generic map ( name => "Block0_complete_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_complete_pipe_read_req(0),
          oack => Block0_complete_pipe_read_ack(0),
          odata => Block0_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_starting_772_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_starting_772_inst_req_0;
      WPIPE_Block0_starting_772_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_starting_772_inst_req_1;
      WPIPE_Block0_starting_772_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= conv_771;
      Block0_starting_write_0_gI: SplitGuardInterface generic map(name => "Block0_starting_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_starting_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_starting", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_starting_pipe_write_req(0),
          oack => Block0_starting_pipe_write_ack(0),
          odata => Block0_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_766_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_766_call_req_0;
      call_stmt_766_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_766_call_req_1;
      call_stmt_766_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_766 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_779_call 
    sendOutput_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_779_call_req_0;
      call_stmt_779_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_779_call_req_1;
      call_stmt_779_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_A is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_A;
architecture zeropad3D_A_arch of zeropad3D_A is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_A_CP_2875_start: Boolean;
  signal zeropad3D_A_CP_2875_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_807_addr_0_ack_0 : boolean;
  signal LOAD_pad_791_load_0_req_1 : boolean;
  signal type_cast_795_inst_req_1 : boolean;
  signal ptr_deref_807_addr_1_ack_1 : boolean;
  signal ptr_deref_807_addr_3_req_1 : boolean;
  signal ptr_deref_1038_store_0_ack_1 : boolean;
  signal LOAD_pad_791_load_0_ack_1 : boolean;
  signal ptr_deref_807_addr_0_req_0 : boolean;
  signal type_cast_795_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_787_inst_req_1 : boolean;
  signal ptr_deref_807_addr_3_ack_0 : boolean;
  signal ptr_deref_807_addr_2_ack_1 : boolean;
  signal ptr_deref_807_addr_2_req_0 : boolean;
  signal ptr_deref_807_addr_3_ack_1 : boolean;
  signal ptr_deref_807_addr_3_req_0 : boolean;
  signal LOAD_pad_791_load_0_ack_0 : boolean;
  signal ptr_deref_807_load_0_ack_0 : boolean;
  signal LOAD_pad_791_load_0_req_0 : boolean;
  signal RPIPE_Block0_starting_787_inst_ack_1 : boolean;
  signal ptr_deref_807_addr_1_ack_0 : boolean;
  signal ptr_deref_807_addr_1_req_1 : boolean;
  signal ptr_deref_807_addr_1_req_0 : boolean;
  signal ptr_deref_807_load_0_req_0 : boolean;
  signal ptr_deref_976_load_3_req_0 : boolean;
  signal ptr_deref_976_addr_2_ack_1 : boolean;
  signal ptr_deref_976_addr_2_req_1 : boolean;
  signal ptr_deref_976_load_3_ack_0 : boolean;
  signal ptr_deref_1038_store_0_ack_0 : boolean;
  signal ptr_deref_976_load_1_ack_1 : boolean;
  signal ptr_deref_976_load_1_req_1 : boolean;
  signal ptr_deref_976_addr_3_req_0 : boolean;
  signal ptr_deref_807_load_1_req_1 : boolean;
  signal ptr_deref_807_addr_2_ack_0 : boolean;
  signal ptr_deref_807_load_2_req_1 : boolean;
  signal ptr_deref_807_load_2_ack_1 : boolean;
  signal ptr_deref_807_load_3_ack_0 : boolean;
  signal RPIPE_Block0_starting_787_inst_req_0 : boolean;
  signal ptr_deref_807_load_0_req_1 : boolean;
  signal RPIPE_Block0_starting_787_inst_ack_0 : boolean;
  signal ptr_deref_807_addr_0_req_1 : boolean;
  signal ptr_deref_807_load_0_ack_1 : boolean;
  signal ptr_deref_807_load_3_req_0 : boolean;
  signal ptr_deref_807_load_1_req_0 : boolean;
  signal type_cast_795_inst_req_0 : boolean;
  signal ptr_deref_976_addr_2_ack_0 : boolean;
  signal ptr_deref_807_load_2_req_0 : boolean;
  signal ptr_deref_807_load_1_ack_1 : boolean;
  signal ptr_deref_807_addr_0_ack_1 : boolean;
  signal type_cast_795_inst_ack_0 : boolean;
  signal ptr_deref_807_load_1_ack_0 : boolean;
  signal ptr_deref_807_addr_2_req_1 : boolean;
  signal ptr_deref_807_load_2_ack_0 : boolean;
  signal addr_of_1113_final_reg_req_0 : boolean;
  signal array_obj_ref_1112_index_offset_req_0 : boolean;
  signal array_obj_ref_1112_index_offset_req_1 : boolean;
  signal addr_of_1113_final_reg_req_1 : boolean;
  signal array_obj_ref_1112_index_offset_ack_0 : boolean;
  signal addr_of_1113_final_reg_ack_0 : boolean;
  signal ptr_deref_1038_store_0_req_0 : boolean;
  signal array_obj_ref_1112_index_offset_ack_1 : boolean;
  signal ptr_deref_976_addr_3_req_1 : boolean;
  signal addr_of_1113_final_reg_ack_1 : boolean;
  signal ptr_deref_976_addr_3_ack_1 : boolean;
  signal ptr_deref_807_load_3_req_1 : boolean;
  signal ptr_deref_807_load_3_ack_1 : boolean;
  signal type_cast_1028_inst_ack_1 : boolean;
  signal type_cast_1028_inst_req_1 : boolean;
  signal type_cast_1106_inst_ack_1 : boolean;
  signal ptr_deref_819_addr_0_req_0 : boolean;
  signal ptr_deref_819_addr_0_ack_0 : boolean;
  signal ptr_deref_976_load_2_ack_0 : boolean;
  signal ptr_deref_819_addr_0_req_1 : boolean;
  signal ptr_deref_819_addr_0_ack_1 : boolean;
  signal type_cast_1106_inst_req_1 : boolean;
  signal type_cast_1028_inst_ack_0 : boolean;
  signal ptr_deref_819_addr_1_req_0 : boolean;
  signal ptr_deref_819_addr_1_ack_0 : boolean;
  signal ptr_deref_976_load_2_req_0 : boolean;
  signal ptr_deref_819_addr_1_req_1 : boolean;
  signal ptr_deref_819_addr_1_ack_1 : boolean;
  signal type_cast_1028_inst_req_0 : boolean;
  signal ptr_deref_819_addr_2_req_0 : boolean;
  signal ptr_deref_819_addr_2_ack_0 : boolean;
  signal ptr_deref_819_addr_2_req_1 : boolean;
  signal addr_of_1035_final_reg_ack_1 : boolean;
  signal ptr_deref_819_addr_2_ack_1 : boolean;
  signal ptr_deref_819_addr_3_req_0 : boolean;
  signal addr_of_1035_final_reg_req_1 : boolean;
  signal ptr_deref_819_addr_3_ack_0 : boolean;
  signal ptr_deref_819_addr_3_req_1 : boolean;
  signal ptr_deref_819_addr_3_ack_1 : boolean;
  signal ptr_deref_976_load_1_ack_0 : boolean;
  signal type_cast_1106_inst_ack_0 : boolean;
  signal type_cast_1106_inst_req_0 : boolean;
  signal ptr_deref_819_load_0_req_0 : boolean;
  signal addr_of_1035_final_reg_ack_0 : boolean;
  signal ptr_deref_819_load_0_ack_0 : boolean;
  signal ptr_deref_819_load_1_req_0 : boolean;
  signal addr_of_1035_final_reg_req_0 : boolean;
  signal ptr_deref_819_load_1_ack_0 : boolean;
  signal ptr_deref_976_load_1_req_0 : boolean;
  signal ptr_deref_819_load_2_req_0 : boolean;
  signal ptr_deref_819_load_2_ack_0 : boolean;
  signal ptr_deref_976_addr_2_req_0 : boolean;
  signal ptr_deref_819_load_3_req_0 : boolean;
  signal ptr_deref_819_load_3_ack_0 : boolean;
  signal ptr_deref_976_load_0_ack_1 : boolean;
  signal ptr_deref_819_load_0_req_1 : boolean;
  signal ptr_deref_819_load_0_ack_1 : boolean;
  signal ptr_deref_819_load_1_req_1 : boolean;
  signal ptr_deref_819_load_1_ack_1 : boolean;
  signal ptr_deref_819_load_2_req_1 : boolean;
  signal ptr_deref_819_load_2_ack_1 : boolean;
  signal ptr_deref_819_load_3_req_1 : boolean;
  signal ptr_deref_819_load_3_ack_1 : boolean;
  signal array_obj_ref_1034_index_offset_ack_1 : boolean;
  signal ptr_deref_976_load_0_ack_0 : boolean;
  signal ptr_deref_976_addr_1_ack_1 : boolean;
  signal ptr_deref_1038_store_0_req_1 : boolean;
  signal ptr_deref_976_addr_3_ack_0 : boolean;
  signal if_stmt_988_branch_ack_0 : boolean;
  signal array_obj_ref_1034_index_offset_req_1 : boolean;
  signal ptr_deref_976_load_0_req_0 : boolean;
  signal ptr_deref_976_addr_1_req_1 : boolean;
  signal if_stmt_988_branch_ack_1 : boolean;
  signal ptr_deref_976_load_0_req_1 : boolean;
  signal ptr_deref_831_load_0_req_0 : boolean;
  signal ptr_deref_831_load_0_ack_0 : boolean;
  signal ptr_deref_831_load_0_req_1 : boolean;
  signal ptr_deref_831_load_0_ack_1 : boolean;
  signal if_stmt_988_branch_req_0 : boolean;
  signal array_obj_ref_1034_index_offset_ack_0 : boolean;
  signal array_obj_ref_1034_index_offset_req_0 : boolean;
  signal ptr_deref_976_load_3_ack_1 : boolean;
  signal ptr_deref_976_load_3_req_1 : boolean;
  signal ptr_deref_976_addr_1_ack_0 : boolean;
  signal ptr_deref_843_load_0_req_0 : boolean;
  signal ptr_deref_843_load_0_ack_0 : boolean;
  signal ptr_deref_976_addr_1_req_0 : boolean;
  signal ptr_deref_843_load_0_req_1 : boolean;
  signal ptr_deref_976_load_2_ack_1 : boolean;
  signal ptr_deref_843_load_0_ack_1 : boolean;
  signal ptr_deref_976_load_2_req_1 : boolean;
  signal ptr_deref_860_addr_0_req_0 : boolean;
  signal ptr_deref_860_addr_0_ack_0 : boolean;
  signal ptr_deref_860_addr_0_req_1 : boolean;
  signal ptr_deref_860_addr_0_ack_1 : boolean;
  signal ptr_deref_860_addr_1_req_0 : boolean;
  signal ptr_deref_860_addr_1_ack_0 : boolean;
  signal ptr_deref_860_addr_1_req_1 : boolean;
  signal ptr_deref_860_addr_1_ack_1 : boolean;
  signal ptr_deref_860_addr_2_req_0 : boolean;
  signal ptr_deref_860_addr_2_ack_0 : boolean;
  signal ptr_deref_860_addr_2_req_1 : boolean;
  signal ptr_deref_860_addr_2_ack_1 : boolean;
  signal ptr_deref_860_addr_3_req_0 : boolean;
  signal ptr_deref_860_addr_3_ack_0 : boolean;
  signal ptr_deref_860_addr_3_req_1 : boolean;
  signal ptr_deref_860_addr_3_ack_1 : boolean;
  signal ptr_deref_860_load_0_req_0 : boolean;
  signal ptr_deref_860_load_0_ack_0 : boolean;
  signal ptr_deref_860_load_1_req_0 : boolean;
  signal ptr_deref_860_load_1_ack_0 : boolean;
  signal ptr_deref_860_load_2_req_0 : boolean;
  signal ptr_deref_860_load_2_ack_0 : boolean;
  signal ptr_deref_860_load_3_req_0 : boolean;
  signal ptr_deref_860_load_3_ack_0 : boolean;
  signal ptr_deref_860_load_0_req_1 : boolean;
  signal ptr_deref_860_load_0_ack_1 : boolean;
  signal ptr_deref_860_load_1_req_1 : boolean;
  signal ptr_deref_860_load_1_ack_1 : boolean;
  signal ptr_deref_860_load_2_req_1 : boolean;
  signal ptr_deref_860_load_2_ack_1 : boolean;
  signal ptr_deref_860_load_3_req_1 : boolean;
  signal ptr_deref_860_load_3_ack_1 : boolean;
  signal if_stmt_879_branch_req_0 : boolean;
  signal if_stmt_879_branch_ack_1 : boolean;
  signal if_stmt_879_branch_ack_0 : boolean;
  signal if_stmt_930_branch_req_0 : boolean;
  signal if_stmt_930_branch_ack_1 : boolean;
  signal if_stmt_930_branch_ack_0 : boolean;
  signal if_stmt_959_branch_req_0 : boolean;
  signal if_stmt_959_branch_ack_1 : boolean;
  signal if_stmt_959_branch_ack_0 : boolean;
  signal ptr_deref_976_addr_0_req_0 : boolean;
  signal ptr_deref_976_addr_0_ack_0 : boolean;
  signal ptr_deref_976_addr_0_req_1 : boolean;
  signal ptr_deref_976_addr_0_ack_1 : boolean;
  signal ptr_deref_1117_load_0_req_0 : boolean;
  signal ptr_deref_1117_load_0_ack_0 : boolean;
  signal ptr_deref_1117_load_0_req_1 : boolean;
  signal ptr_deref_1117_load_0_ack_1 : boolean;
  signal type_cast_1131_inst_req_0 : boolean;
  signal type_cast_1131_inst_ack_0 : boolean;
  signal type_cast_1131_inst_req_1 : boolean;
  signal type_cast_1131_inst_ack_1 : boolean;
  signal array_obj_ref_1137_index_offset_req_0 : boolean;
  signal array_obj_ref_1137_index_offset_ack_0 : boolean;
  signal array_obj_ref_1137_index_offset_req_1 : boolean;
  signal array_obj_ref_1137_index_offset_ack_1 : boolean;
  signal addr_of_1138_final_reg_req_0 : boolean;
  signal addr_of_1138_final_reg_ack_0 : boolean;
  signal addr_of_1138_final_reg_req_1 : boolean;
  signal addr_of_1138_final_reg_ack_1 : boolean;
  signal ptr_deref_1141_store_0_req_0 : boolean;
  signal ptr_deref_1141_store_0_ack_0 : boolean;
  signal ptr_deref_1141_store_0_req_1 : boolean;
  signal ptr_deref_1141_store_0_ack_1 : boolean;
  signal if_stmt_1159_branch_req_0 : boolean;
  signal if_stmt_1159_branch_ack_1 : boolean;
  signal if_stmt_1159_branch_ack_0 : boolean;
  signal ptr_deref_1182_addr_0_req_0 : boolean;
  signal ptr_deref_1182_addr_0_ack_0 : boolean;
  signal ptr_deref_1182_addr_0_req_1 : boolean;
  signal ptr_deref_1182_addr_0_ack_1 : boolean;
  signal ptr_deref_1182_addr_1_req_0 : boolean;
  signal ptr_deref_1182_addr_1_ack_0 : boolean;
  signal ptr_deref_1182_addr_1_req_1 : boolean;
  signal ptr_deref_1182_addr_1_ack_1 : boolean;
  signal ptr_deref_1182_addr_2_req_0 : boolean;
  signal ptr_deref_1182_addr_2_ack_0 : boolean;
  signal ptr_deref_1182_addr_2_req_1 : boolean;
  signal ptr_deref_1182_addr_2_ack_1 : boolean;
  signal ptr_deref_1182_addr_3_req_0 : boolean;
  signal ptr_deref_1182_addr_3_ack_0 : boolean;
  signal ptr_deref_1182_addr_3_req_1 : boolean;
  signal ptr_deref_1182_addr_3_ack_1 : boolean;
  signal ptr_deref_1182_load_0_req_0 : boolean;
  signal ptr_deref_1182_load_0_ack_0 : boolean;
  signal ptr_deref_1182_load_1_req_0 : boolean;
  signal ptr_deref_1182_load_1_ack_0 : boolean;
  signal ptr_deref_1182_load_2_req_0 : boolean;
  signal ptr_deref_1182_load_2_ack_0 : boolean;
  signal ptr_deref_1182_load_3_req_0 : boolean;
  signal ptr_deref_1182_load_3_ack_0 : boolean;
  signal ptr_deref_1182_load_0_req_1 : boolean;
  signal ptr_deref_1182_load_0_ack_1 : boolean;
  signal ptr_deref_1182_load_1_req_1 : boolean;
  signal ptr_deref_1182_load_1_ack_1 : boolean;
  signal ptr_deref_1182_load_2_req_1 : boolean;
  signal ptr_deref_1182_load_2_ack_1 : boolean;
  signal ptr_deref_1182_load_3_req_1 : boolean;
  signal ptr_deref_1182_load_3_ack_1 : boolean;
  signal type_cast_1196_inst_req_0 : boolean;
  signal type_cast_1196_inst_ack_0 : boolean;
  signal type_cast_1196_inst_req_1 : boolean;
  signal type_cast_1196_inst_ack_1 : boolean;
  signal if_stmt_1203_branch_req_0 : boolean;
  signal if_stmt_1203_branch_ack_1 : boolean;
  signal if_stmt_1203_branch_ack_0 : boolean;
  signal ptr_deref_1250_addr_0_req_0 : boolean;
  signal ptr_deref_1250_addr_0_ack_0 : boolean;
  signal ptr_deref_1250_addr_0_req_1 : boolean;
  signal ptr_deref_1250_addr_0_ack_1 : boolean;
  signal ptr_deref_1250_addr_1_req_0 : boolean;
  signal ptr_deref_1250_addr_1_ack_0 : boolean;
  signal ptr_deref_1250_addr_1_req_1 : boolean;
  signal ptr_deref_1250_addr_1_ack_1 : boolean;
  signal ptr_deref_1250_addr_2_req_0 : boolean;
  signal ptr_deref_1250_addr_2_ack_0 : boolean;
  signal ptr_deref_1250_addr_2_req_1 : boolean;
  signal ptr_deref_1250_addr_2_ack_1 : boolean;
  signal ptr_deref_1250_addr_3_req_0 : boolean;
  signal ptr_deref_1250_addr_3_ack_0 : boolean;
  signal ptr_deref_1250_addr_3_req_1 : boolean;
  signal ptr_deref_1250_addr_3_ack_1 : boolean;
  signal ptr_deref_1250_load_0_req_0 : boolean;
  signal ptr_deref_1250_load_0_ack_0 : boolean;
  signal ptr_deref_1250_load_1_req_0 : boolean;
  signal ptr_deref_1250_load_1_ack_0 : boolean;
  signal ptr_deref_1250_load_2_req_0 : boolean;
  signal ptr_deref_1250_load_2_ack_0 : boolean;
  signal ptr_deref_1250_load_3_req_0 : boolean;
  signal ptr_deref_1250_load_3_ack_0 : boolean;
  signal ptr_deref_1250_load_0_req_1 : boolean;
  signal ptr_deref_1250_load_0_ack_1 : boolean;
  signal ptr_deref_1250_load_1_req_1 : boolean;
  signal ptr_deref_1250_load_1_ack_1 : boolean;
  signal ptr_deref_1250_load_2_req_1 : boolean;
  signal ptr_deref_1250_load_2_ack_1 : boolean;
  signal ptr_deref_1250_load_3_req_1 : boolean;
  signal ptr_deref_1250_load_3_ack_1 : boolean;
  signal if_stmt_1262_branch_req_0 : boolean;
  signal if_stmt_1262_branch_ack_1 : boolean;
  signal if_stmt_1262_branch_ack_0 : boolean;
  signal WPIPE_Block0_complete_1272_inst_req_0 : boolean;
  signal WPIPE_Block0_complete_1272_inst_ack_0 : boolean;
  signal WPIPE_Block0_complete_1272_inst_req_1 : boolean;
  signal WPIPE_Block0_complete_1272_inst_ack_1 : boolean;
  signal type_cast_897_inst_req_0 : boolean;
  signal type_cast_897_inst_ack_0 : boolean;
  signal type_cast_897_inst_req_1 : boolean;
  signal type_cast_897_inst_ack_1 : boolean;
  signal phi_stmt_894_req_0 : boolean;
  signal phi_stmt_900_req_0 : boolean;
  signal phi_stmt_907_req_0 : boolean;
  signal phi_stmt_914_req_0 : boolean;
  signal type_cast_899_inst_req_0 : boolean;
  signal type_cast_899_inst_ack_0 : boolean;
  signal type_cast_899_inst_req_1 : boolean;
  signal type_cast_899_inst_ack_1 : boolean;
  signal phi_stmt_894_req_1 : boolean;
  signal type_cast_906_inst_req_0 : boolean;
  signal type_cast_906_inst_ack_0 : boolean;
  signal type_cast_906_inst_req_1 : boolean;
  signal type_cast_906_inst_ack_1 : boolean;
  signal phi_stmt_900_req_1 : boolean;
  signal type_cast_913_inst_req_0 : boolean;
  signal type_cast_913_inst_ack_0 : boolean;
  signal type_cast_913_inst_req_1 : boolean;
  signal type_cast_913_inst_ack_1 : boolean;
  signal phi_stmt_907_req_1 : boolean;
  signal type_cast_920_inst_req_0 : boolean;
  signal type_cast_920_inst_ack_0 : boolean;
  signal type_cast_920_inst_req_1 : boolean;
  signal type_cast_920_inst_ack_1 : boolean;
  signal phi_stmt_914_req_1 : boolean;
  signal phi_stmt_894_ack_0 : boolean;
  signal phi_stmt_900_ack_0 : boolean;
  signal phi_stmt_907_ack_0 : boolean;
  signal phi_stmt_914_ack_0 : boolean;
  signal type_cast_1220_inst_req_0 : boolean;
  signal type_cast_1220_inst_ack_0 : boolean;
  signal type_cast_1220_inst_req_1 : boolean;
  signal type_cast_1220_inst_ack_1 : boolean;
  signal phi_stmt_1212_req_2 : boolean;
  signal type_cast_1230_inst_req_0 : boolean;
  signal type_cast_1230_inst_ack_0 : boolean;
  signal type_cast_1230_inst_req_1 : boolean;
  signal type_cast_1230_inst_ack_1 : boolean;
  signal phi_stmt_1221_req_2 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal phi_stmt_1231_req_2 : boolean;
  signal type_cast_1218_inst_req_0 : boolean;
  signal type_cast_1218_inst_ack_0 : boolean;
  signal type_cast_1218_inst_req_1 : boolean;
  signal type_cast_1218_inst_ack_1 : boolean;
  signal phi_stmt_1212_req_1 : boolean;
  signal phi_stmt_1221_req_1 : boolean;
  signal type_cast_1236_inst_req_0 : boolean;
  signal type_cast_1236_inst_ack_0 : boolean;
  signal type_cast_1236_inst_req_1 : boolean;
  signal type_cast_1236_inst_ack_1 : boolean;
  signal phi_stmt_1231_req_1 : boolean;
  signal phi_stmt_1212_req_0 : boolean;
  signal phi_stmt_1221_req_0 : boolean;
  signal type_cast_1234_inst_req_0 : boolean;
  signal type_cast_1234_inst_ack_0 : boolean;
  signal type_cast_1234_inst_req_1 : boolean;
  signal type_cast_1234_inst_ack_1 : boolean;
  signal phi_stmt_1231_req_0 : boolean;
  signal phi_stmt_1212_ack_0 : boolean;
  signal phi_stmt_1221_ack_0 : boolean;
  signal phi_stmt_1231_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_A_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_A_CP_2875_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_A_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2875_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2875_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_2875_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_A_CP_2875: Block -- control-path 
    signal zeropad3D_A_CP_2875_elements: BooleanArray(243 downto 0);
    -- 
  begin -- 
    zeropad3D_A_CP_2875_elements(0) <= zeropad3D_A_CP_2875_start;
    zeropad3D_A_CP_2875_symbol <= zeropad3D_A_CP_2875_elements(185);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_785/assign_stmt_788__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_785/assign_stmt_788/$entry
      -- CP-element group 0: 	 branch_block_stmt_785/branch_block_stmt_785__entry__
      -- CP-element group 0: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_785/$entry
      -- CP-element group 0: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_Sample/rr
      -- 
    rr_2957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(0), ack => RPIPE_Block0_starting_787_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_update_start_
      -- CP-element group 1: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_Update/$entry
      -- 
    ra_2958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_787_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(1)); -- 
    cr_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(1), ack => RPIPE_Block0_starting_787_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	35 
    -- CP-element group 2: 	36 
    -- CP-element group 2: 	37 
    -- CP-element group 2: 	33 
    -- CP-element group 2: 	34 
    -- CP-element group 2: 	71 
    -- CP-element group 2: 	72 
    -- CP-element group 2: 	31 
    -- CP-element group 2: 	32 
    -- CP-element group 2: 	38 
    -- CP-element group 2: 	69 
    -- CP-element group 2: 	70 
    -- CP-element group 2: 	44 
    -- CP-element group 2: 	45 
    -- CP-element group 2: 	46 
    -- CP-element group 2: 	47 
    -- CP-element group 2: 	49 
    -- CP-element group 2: 	50 
    -- CP-element group 2: 	51 
    -- CP-element group 2: 	52 
    -- CP-element group 2: 	53 
    -- CP-element group 2: 	56 
    -- CP-element group 2: 	57 
    -- CP-element group 2: 	58 
    -- CP-element group 2: 	59 
    -- CP-element group 2: 	60 
    -- CP-element group 2: 	61 
    -- CP-element group 2: 	62 
    -- CP-element group 2: 	63 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2:  members (194) 
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_0_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_1_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_3_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_0_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_788/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_2_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_788__exit__
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_update_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_update_start
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_2_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_3_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_3_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_sample_start
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_1_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_1_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878__entry__
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_update_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_0_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_1/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_2/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_3_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_0_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_2/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_2_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_788/RPIPE_Block0_starting_787_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_1/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_1_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_2_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_update_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_3/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_3/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_update_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_sample_start
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_update_start
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_0_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_0_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_0_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_0_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_1_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_1_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_1_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_1_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_2_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_2_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_2_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_2_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_3_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_3_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_3_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_3_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_1/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_1/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_2/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_2/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_3/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_3/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_update_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_update_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_update_start_
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_sample_start
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_update_start
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_0_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_0_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_0_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_0_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_1_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_1_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_1_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_1_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_2_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_2_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_2_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_2_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_3_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_3_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_3_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_3_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_1/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_1/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_2/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_2/cr
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_3/$entry
      -- CP-element group 2: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_3/cr
      -- 
    ca_2963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_787_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(2)); -- 
    cr_2993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => LOAD_pad_791_load_0_req_1); -- 
    cr_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => type_cast_795_inst_req_1); -- 
    cr_3074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_addr_3_req_1); -- 
    rr_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_addr_0_req_0); -- 
    rr_3059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_addr_2_req_0); -- 
    rr_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_addr_3_req_0); -- 
    rr_2982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => LOAD_pad_791_load_0_req_0); -- 
    cr_3054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_addr_1_req_1); -- 
    rr_3049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_addr_1_req_0); -- 
    cr_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_load_1_req_1); -- 
    cr_3121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_load_2_req_1); -- 
    cr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_load_0_req_1); -- 
    cr_3044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_addr_0_req_1); -- 
    cr_3064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_addr_2_req_1); -- 
    cr_3126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_807_load_3_req_1); -- 
    rr_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_addr_0_req_0); -- 
    cr_3163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_addr_0_req_1); -- 
    rr_3168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_addr_1_req_0); -- 
    cr_3173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_addr_1_req_1); -- 
    rr_3178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_addr_2_req_0); -- 
    cr_3183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_addr_2_req_1); -- 
    rr_3188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_addr_3_req_0); -- 
    cr_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_addr_3_req_1); -- 
    cr_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_load_0_req_1); -- 
    cr_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_load_1_req_1); -- 
    cr_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_load_2_req_1); -- 
    cr_3245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_819_load_3_req_1); -- 
    rr_3284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_831_load_0_req_0); -- 
    cr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_831_load_0_req_1); -- 
    rr_3334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_843_load_0_req_0); -- 
    cr_3345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_843_load_0_req_1); -- 
    rr_3377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_addr_0_req_0); -- 
    cr_3382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_addr_0_req_1); -- 
    rr_3387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_addr_1_req_0); -- 
    cr_3392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_addr_1_req_1); -- 
    rr_3397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_addr_2_req_0); -- 
    cr_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_addr_2_req_1); -- 
    rr_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_addr_3_req_0); -- 
    cr_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_addr_3_req_1); -- 
    cr_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_load_0_req_1); -- 
    cr_3454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_load_1_req_1); -- 
    cr_3459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_load_2_req_1); -- 
    cr_3464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(2), ack => ptr_deref_860_load_3_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Sample/word_access_start/word_0/ra
      -- 
    ra_2983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_791_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/LOAD_pad_791_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/LOAD_pad_791_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/LOAD_pad_791_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/LOAD_pad_791_Update/LOAD_pad_791_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_Sample/rr
      -- 
    ca_2994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_791_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(4)); -- 
    rr_3007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(4), ack => type_cast_795_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_Sample/ra
      -- 
    ra_3008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_795_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	74 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/type_cast_795_Update/$exit
      -- 
    ca_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_795_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(6)); -- 
    -- CP-element group 7:  join  fork  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	9 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	18 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	21 
    -- CP-element group 7:  members (11) 
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_1/$entry
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_0/rr
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_3/rr
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_1/rr
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_2/rr
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_2/$entry
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_3/$entry
      -- CP-element group 7: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/$entry
      -- 
    rr_3085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(7), ack => ptr_deref_807_load_0_req_0); -- 
    rr_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(7), ack => ptr_deref_807_load_1_req_0); -- 
    rr_3095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(7), ack => ptr_deref_807_load_2_req_0); -- 
    rr_3100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(7), ack => ptr_deref_807_load_3_req_0); -- 
    zeropad3D_A_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_A_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(2) & zeropad3D_A_CP_2875_elements(9);
      gj_zeropad3D_A_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  transition  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: 	12 
    -- CP-element group 8: 	14 
    -- CP-element group 8: 	16 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	74 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_sample_complete
      -- 
    zeropad3D_A_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_A_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(10) & zeropad3D_A_CP_2875_elements(12) & zeropad3D_A_CP_2875_elements(14) & zeropad3D_A_CP_2875_elements(16);
      gj_zeropad3D_A_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	17 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_update_complete
      -- CP-element group 9: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_address_calculated
      -- 
    zeropad3D_A_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_A_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(11) & zeropad3D_A_CP_2875_elements(13) & zeropad3D_A_CP_2875_elements(15) & zeropad3D_A_CP_2875_elements(17);
      gj_zeropad3D_A_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_0_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_0_Sample/$exit
      -- 
    ra_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_addr_0_ack_0, ack => zeropad3D_A_CP_2875_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_0_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_0_Update/ca
      -- 
    ca_3045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_addr_0_ack_1, ack => zeropad3D_A_CP_2875_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_1_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_1_Sample/$exit
      -- 
    ra_3050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_addr_1_ack_0, ack => zeropad3D_A_CP_2875_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	9 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_1_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_1_Update/$exit
      -- 
    ca_3055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_addr_1_ack_1, ack => zeropad3D_A_CP_2875_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	8 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_2_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_2_Sample/ra
      -- 
    ra_3060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_addr_2_ack_0, ack => zeropad3D_A_CP_2875_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	9 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_2_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_2_Update/$exit
      -- 
    ca_3065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_addr_2_ack_1, ack => zeropad3D_A_CP_2875_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	8 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_3_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_3_Sample/$exit
      -- 
    ra_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_addr_3_ack_0, ack => zeropad3D_A_CP_2875_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	9 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_3_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_word_addrgen_3_Update/ca
      -- 
    ca_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_addr_3_ack_1, ack => zeropad3D_A_CP_2875_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	7 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_0/ra
      -- CP-element group 18: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_0/$exit
      -- 
    ra_3086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_1/$exit
      -- CP-element group 19: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_1/ra
      -- 
    ra_3091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_load_1_ack_0, ack => zeropad3D_A_CP_2875_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_2/$exit
      -- CP-element group 20: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_2/ra
      -- 
    ra_3096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_load_2_ack_0, ack => zeropad3D_A_CP_2875_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_3/ra
      -- CP-element group 21: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/word_3/$exit
      -- 
    ra_3101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_load_3_ack_0, ack => zeropad3D_A_CP_2875_elements(21)); -- 
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/word_access_start/$exit
      -- CP-element group 22: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Sample/$exit
      -- 
    zeropad3D_A_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(18) & zeropad3D_A_CP_2875_elements(19) & zeropad3D_A_CP_2875_elements(20) & zeropad3D_A_CP_2875_elements(21);
      gj_zeropad3D_A_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	27 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_0/ca
      -- CP-element group 23: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_0/$exit
      -- 
    ca_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	27 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_1/$exit
      -- CP-element group 24: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_1/ca
      -- 
    ca_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_load_1_ack_1, ack => zeropad3D_A_CP_2875_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_2/ca
      -- CP-element group 25: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_2/$exit
      -- 
    ca_3122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_load_2_ack_1, ack => zeropad3D_A_CP_2875_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_3/$exit
      -- CP-element group 26: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/word_3/ca
      -- 
    ca_3127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_807_load_3_ack_1, ack => zeropad3D_A_CP_2875_elements(26)); -- 
    -- CP-element group 27:  join  transition  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: 	24 
    -- CP-element group 27: 	25 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	74 
    -- CP-element group 27:  members (7) 
      -- CP-element group 27: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/word_access_complete/$exit
      -- CP-element group 27: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/ptr_deref_807_Merge/$entry
      -- CP-element group 27: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/ptr_deref_807_Merge/$exit
      -- CP-element group 27: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/ptr_deref_807_Merge/merge_req
      -- CP-element group 27: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_807_Update/ptr_deref_807_Merge/merge_ack
      -- 
    zeropad3D_A_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(23) & zeropad3D_A_CP_2875_elements(24) & zeropad3D_A_CP_2875_elements(25) & zeropad3D_A_CP_2875_elements(26);
      gj_zeropad3D_A_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	39 
    -- CP-element group 28: 	40 
    -- CP-element group 28: 	41 
    -- CP-element group 28: 	42 
    -- CP-element group 28:  members (11) 
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/$entry
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_0/$entry
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_0/rr
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_1/$entry
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_1/rr
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_2/$entry
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_2/rr
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_3/$entry
      -- CP-element group 28: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_3/rr
      -- 
    rr_3204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(28), ack => ptr_deref_819_load_0_req_0); -- 
    rr_3209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(28), ack => ptr_deref_819_load_1_req_0); -- 
    rr_3214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(28), ack => ptr_deref_819_load_2_req_0); -- 
    rr_3219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(28), ack => ptr_deref_819_load_3_req_0); -- 
    zeropad3D_A_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(30) & zeropad3D_A_CP_2875_elements(2);
      gj_zeropad3D_A_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	35 
    -- CP-element group 29: 	37 
    -- CP-element group 29: 	33 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	74 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_sample_complete
      -- 
    zeropad3D_A_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(35) & zeropad3D_A_CP_2875_elements(37) & zeropad3D_A_CP_2875_elements(33) & zeropad3D_A_CP_2875_elements(31);
      gj_zeropad3D_A_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	36 
    -- CP-element group 30: 	34 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	38 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_address_calculated
      -- CP-element group 30: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_update_complete
      -- 
    zeropad3D_A_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(36) & zeropad3D_A_CP_2875_elements(34) & zeropad3D_A_CP_2875_elements(32) & zeropad3D_A_CP_2875_elements(38);
      gj_zeropad3D_A_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	2 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_0_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_0_Sample/ra
      -- 
    ra_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_addr_0_ack_0, ack => zeropad3D_A_CP_2875_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_0_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_0_Update/ca
      -- 
    ca_3164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_addr_0_ack_1, ack => zeropad3D_A_CP_2875_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	2 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	29 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_1_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_1_Sample/ra
      -- 
    ra_3169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_addr_1_ack_0, ack => zeropad3D_A_CP_2875_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	2 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	30 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_1_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_1_Update/ca
      -- 
    ca_3174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_addr_1_ack_1, ack => zeropad3D_A_CP_2875_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	2 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	29 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_2_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_2_Sample/ra
      -- 
    ra_3179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_addr_2_ack_0, ack => zeropad3D_A_CP_2875_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	2 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	30 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_2_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_2_Update/ca
      -- 
    ca_3184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_addr_2_ack_1, ack => zeropad3D_A_CP_2875_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	2 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	29 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_3_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_3_Sample/ra
      -- 
    ra_3189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_addr_3_ack_0, ack => zeropad3D_A_CP_2875_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	2 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	30 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_3_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_word_addrgen_3_Update/ca
      -- 
    ca_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_addr_3_ack_1, ack => zeropad3D_A_CP_2875_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	28 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	43 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_0/ra
      -- 
    ra_3205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	28 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_1/ra
      -- 
    ra_3210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_load_1_ack_0, ack => zeropad3D_A_CP_2875_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	28 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_2/$exit
      -- CP-element group 41: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_2/ra
      -- 
    ra_3215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_load_2_ack_0, ack => zeropad3D_A_CP_2875_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	28 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_3/$exit
      -- CP-element group 42: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/word_3/ra
      -- 
    ra_3220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_load_3_ack_0, ack => zeropad3D_A_CP_2875_elements(42)); -- 
    -- CP-element group 43:  join  transition  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	39 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	41 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Sample/word_access_start/$exit
      -- 
    zeropad3D_A_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(39) & zeropad3D_A_CP_2875_elements(40) & zeropad3D_A_CP_2875_elements(41) & zeropad3D_A_CP_2875_elements(42);
      gj_zeropad3D_A_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	2 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	48 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_0/ca
      -- 
    ca_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	2 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	48 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_1/ca
      -- 
    ca_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_load_1_ack_1, ack => zeropad3D_A_CP_2875_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	2 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_2/$exit
      -- CP-element group 46: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_2/ca
      -- 
    ca_3241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_load_2_ack_1, ack => zeropad3D_A_CP_2875_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	2 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_3/$exit
      -- CP-element group 47: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/word_3/ca
      -- 
    ca_3246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_819_load_3_ack_1, ack => zeropad3D_A_CP_2875_elements(47)); -- 
    -- CP-element group 48:  join  transition  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	44 
    -- CP-element group 48: 	45 
    -- CP-element group 48: 	46 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (7) 
      -- CP-element group 48: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/ptr_deref_819_Merge/$entry
      -- CP-element group 48: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/ptr_deref_819_Merge/$exit
      -- CP-element group 48: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/ptr_deref_819_Merge/merge_req
      -- CP-element group 48: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_819_Update/ptr_deref_819_Merge/merge_ack
      -- 
    zeropad3D_A_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(44) & zeropad3D_A_CP_2875_elements(45) & zeropad3D_A_CP_2875_elements(46) & zeropad3D_A_CP_2875_elements(47);
      gj_zeropad3D_A_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	2 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Sample/word_access_start/word_0/ra
      -- 
    ra_3285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_831_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	2 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	74 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/word_access_complete/word_0/ca
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/ptr_deref_831_Merge/$entry
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/ptr_deref_831_Merge/$exit
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/ptr_deref_831_Merge/merge_req
      -- CP-element group 50: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_831_Update/ptr_deref_831_Merge/merge_ack
      -- 
    ca_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_831_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	2 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Sample/word_access_start/word_0/ra
      -- 
    ra_3335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_843_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	2 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (9) 
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/word_access_complete/word_0/ca
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/ptr_deref_843_Merge/$entry
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/ptr_deref_843_Merge/$exit
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/ptr_deref_843_Merge/merge_req
      -- CP-element group 52: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_843_Update/ptr_deref_843_Merge/merge_ack
      -- 
    ca_3346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_843_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	2 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	66 
    -- CP-element group 53: 	67 
    -- CP-element group 53: 	64 
    -- CP-element group 53: 	65 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_0/rr
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_1/$entry
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_1/rr
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_2/$entry
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_2/rr
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_3/$entry
      -- CP-element group 53: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_3/rr
      -- 
    rr_3433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(53), ack => ptr_deref_860_load_2_req_0); -- 
    rr_3438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(53), ack => ptr_deref_860_load_3_req_0); -- 
    rr_3423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(53), ack => ptr_deref_860_load_0_req_0); -- 
    rr_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(53), ack => ptr_deref_860_load_1_req_0); -- 
    zeropad3D_A_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(55) & zeropad3D_A_CP_2875_elements(2);
      gj_zeropad3D_A_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: 	58 
    -- CP-element group 54: 	60 
    -- CP-element group 54: 	62 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	74 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_sample_complete
      -- 
    zeropad3D_A_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(56) & zeropad3D_A_CP_2875_elements(58) & zeropad3D_A_CP_2875_elements(60) & zeropad3D_A_CP_2875_elements(62);
      gj_zeropad3D_A_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	57 
    -- CP-element group 55: 	59 
    -- CP-element group 55: 	61 
    -- CP-element group 55: 	63 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_update_complete
      -- 
    zeropad3D_A_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(57) & zeropad3D_A_CP_2875_elements(59) & zeropad3D_A_CP_2875_elements(61) & zeropad3D_A_CP_2875_elements(63);
      gj_zeropad3D_A_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	2 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_0_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_0_Sample/ra
      -- 
    ra_3378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_addr_0_ack_0, ack => zeropad3D_A_CP_2875_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	2 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	55 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_0_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_0_Update/ca
      -- 
    ca_3383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_addr_0_ack_1, ack => zeropad3D_A_CP_2875_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	2 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	54 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_1_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_1_Sample/ra
      -- 
    ra_3388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_addr_1_ack_0, ack => zeropad3D_A_CP_2875_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	55 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_1_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_1_Update/ca
      -- 
    ca_3393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_addr_1_ack_1, ack => zeropad3D_A_CP_2875_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	2 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	54 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_2_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_2_Sample/ra
      -- 
    ra_3398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_addr_2_ack_0, ack => zeropad3D_A_CP_2875_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	2 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	55 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_2_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_2_Update/ca
      -- 
    ca_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_addr_2_ack_1, ack => zeropad3D_A_CP_2875_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	2 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	54 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_3_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_3_Sample/ra
      -- 
    ra_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_addr_3_ack_0, ack => zeropad3D_A_CP_2875_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	2 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	55 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_3_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_word_addrgen_3_Update/ca
      -- 
    ca_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_addr_3_ack_1, ack => zeropad3D_A_CP_2875_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	53 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	68 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_0/ra
      -- 
    ra_3424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	53 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_1/ra
      -- 
    ra_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_1_ack_0, ack => zeropad3D_A_CP_2875_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	53 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_2/$exit
      -- CP-element group 66: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_2/ra
      -- 
    ra_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_2_ack_0, ack => zeropad3D_A_CP_2875_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	53 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_3/$exit
      -- CP-element group 67: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/word_3/ra
      -- 
    ra_3439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_3_ack_0, ack => zeropad3D_A_CP_2875_elements(67)); -- 
    -- CP-element group 68:  join  transition  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	67 
    -- CP-element group 68: 	64 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Sample/word_access_start/$exit
      -- 
    zeropad3D_A_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(66) & zeropad3D_A_CP_2875_elements(67) & zeropad3D_A_CP_2875_elements(64) & zeropad3D_A_CP_2875_elements(65);
      gj_zeropad3D_A_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	2 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	73 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_0/ca
      -- 
    ca_3450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	2 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	73 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_1/$exit
      -- CP-element group 70: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_1/ca
      -- 
    ca_3455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_1_ack_1, ack => zeropad3D_A_CP_2875_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	2 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_2/$exit
      -- CP-element group 71: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_2/ca
      -- 
    ca_3460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_2_ack_1, ack => zeropad3D_A_CP_2875_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	2 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_3/$exit
      -- CP-element group 72: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/word_3/ca
      -- 
    ca_3465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_860_load_3_ack_1, ack => zeropad3D_A_CP_2875_elements(72)); -- 
    -- CP-element group 73:  join  transition  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: 	69 
    -- CP-element group 73: 	70 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (7) 
      -- CP-element group 73: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/word_access_complete/$exit
      -- CP-element group 73: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/ptr_deref_860_Merge/$entry
      -- CP-element group 73: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/ptr_deref_860_Merge/$exit
      -- CP-element group 73: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/ptr_deref_860_Merge/merge_req
      -- CP-element group 73: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/ptr_deref_860_Update/ptr_deref_860_Merge/merge_ack
      -- 
    zeropad3D_A_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(71) & zeropad3D_A_CP_2875_elements(72) & zeropad3D_A_CP_2875_elements(69) & zeropad3D_A_CP_2875_elements(70);
      gj_zeropad3D_A_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	29 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	50 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	54 
    -- CP-element group 74: 	6 
    -- CP-element group 74: 	8 
    -- CP-element group 74: 	27 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878/$exit
      -- CP-element group 74: 	 branch_block_stmt_785/assign_stmt_792_to_assign_stmt_878__exit__
      -- CP-element group 74: 	 branch_block_stmt_785/if_stmt_879__entry__
      -- CP-element group 74: 	 branch_block_stmt_785/if_stmt_879_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_785/if_stmt_879_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_785/if_stmt_879_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_785/if_stmt_879_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_785/R_cmp123_880_place
      -- CP-element group 74: 	 branch_block_stmt_785/if_stmt_879_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_785/if_stmt_879_else_link/$entry
      -- 
    branch_req_3478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(74), ack => if_stmt_879_branch_req_0); -- 
    zeropad3D_A_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(73) & zeropad3D_A_CP_2875_elements(29) & zeropad3D_A_CP_2875_elements(48) & zeropad3D_A_CP_2875_elements(50) & zeropad3D_A_CP_2875_elements(52) & zeropad3D_A_CP_2875_elements(54) & zeropad3D_A_CP_2875_elements(6) & zeropad3D_A_CP_2875_elements(8) & zeropad3D_A_CP_2875_elements(27);
      gj_zeropad3D_A_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  place  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	243 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_785/if_stmt_879_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_785/if_stmt_879_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_785/entry_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_785/entry_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_785/entry_whilex_xend_PhiReq/$entry
      -- 
    if_choice_transition_3483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_879_branch_ack_1, ack => zeropad3D_A_CP_2875_elements(75)); -- 
    -- CP-element group 76:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	190 
    -- CP-element group 76: 	191 
    -- CP-element group 76: 	189 
    -- CP-element group 76: 	186 
    -- CP-element group 76: 	187 
    -- CP-element group 76:  members (30) 
      -- CP-element group 76: 	 branch_block_stmt_785/merge_stmt_885__exit__
      -- CP-element group 76: 	 branch_block_stmt_785/assign_stmt_891__entry__
      -- CP-element group 76: 	 branch_block_stmt_785/assign_stmt_891__exit__
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody
      -- CP-element group 76: 	 branch_block_stmt_785/if_stmt_879_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_785/if_stmt_879_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_785/entry_bbx_xnph
      -- CP-element group 76: 	 branch_block_stmt_785/assign_stmt_891/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/assign_stmt_891/$exit
      -- CP-element group 76: 	 branch_block_stmt_785/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 76: 	 branch_block_stmt_785/merge_stmt_885_PhiReqMerge
      -- CP-element group 76: 	 branch_block_stmt_785/merge_stmt_885_PhiAck/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/merge_stmt_885_PhiAck/$exit
      -- CP-element group 76: 	 branch_block_stmt_785/merge_stmt_885_PhiAck/dummy
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_900/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_907/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_914/$entry
      -- CP-element group 76: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/$entry
      -- 
    else_choice_transition_3487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_879_branch_ack_0, ack => zeropad3D_A_CP_2875_elements(76)); -- 
    rr_4379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(76), ack => type_cast_897_inst_req_0); -- 
    cr_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(76), ack => type_cast_897_inst_req_1); -- 
    -- CP-element group 77:  merge  branch  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	211 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	80 
    -- CP-element group 77:  members (22) 
      -- CP-element group 77: 	 branch_block_stmt_785/assign_stmt_941_to_assign_stmt_958__entry__
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_959__entry__
      -- CP-element group 77: 	 branch_block_stmt_785/merge_stmt_936__exit__
      -- CP-element group 77: 	 branch_block_stmt_785/assign_stmt_941_to_assign_stmt_958__exit__
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_930_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_930_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_785/whilex_xbody_lorx_xlhsx_xfalse
      -- CP-element group 77: 	 branch_block_stmt_785/assign_stmt_941_to_assign_stmt_958/$entry
      -- CP-element group 77: 	 branch_block_stmt_785/assign_stmt_941_to_assign_stmt_958/$exit
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_959_dead_link/$entry
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_959_eval_test/$entry
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_959_eval_test/$exit
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_959_eval_test/branch_req
      -- CP-element group 77: 	 branch_block_stmt_785/R_orx_xcond_960_place
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_959_if_link/$entry
      -- CP-element group 77: 	 branch_block_stmt_785/if_stmt_959_else_link/$entry
      -- CP-element group 77: 	 branch_block_stmt_785/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_785/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_785/merge_stmt_936_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_785/merge_stmt_936_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_785/merge_stmt_936_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_785/merge_stmt_936_PhiAck/dummy
      -- 
    if_choice_transition_3508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_930_branch_ack_1, ack => zeropad3D_A_CP_2875_elements(77)); -- 
    branch_req_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(77), ack => if_stmt_959_branch_req_0); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	211 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	212 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_785/if_stmt_930_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_785/if_stmt_930_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_785/whilex_xbody_ifx_xthen
      -- CP-element group 78: 	 branch_block_stmt_785/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_785/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_930_branch_ack_0, ack => zeropad3D_A_CP_2875_elements(78)); -- 
    -- CP-element group 79:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	99 
    -- CP-element group 79: 	100 
    -- CP-element group 79: 	81 
    -- CP-element group 79: 	84 
    -- CP-element group 79: 	85 
    -- CP-element group 79: 	86 
    -- CP-element group 79: 	87 
    -- CP-element group 79: 	88 
    -- CP-element group 79: 	89 
    -- CP-element group 79: 	90 
    -- CP-element group 79: 	91 
    -- CP-element group 79: 	97 
    -- CP-element group 79: 	98 
    -- CP-element group 79:  members (52) 
      -- CP-element group 79: 	 branch_block_stmt_785/merge_stmt_965__exit__
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_2_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_2_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_1/cr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_3_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_3_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987__entry__
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_1_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_2/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_3_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_3_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_1/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_2_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_2_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_1_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_0/cr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_0/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_1_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_3/cr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_3/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_1_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_2/cr
      -- CP-element group 79: 	 branch_block_stmt_785/if_stmt_959_if_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_785/if_stmt_959_if_link/if_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_785/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse43
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_update_start_
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_address_calculated
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_root_address_calculated
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_address_resized
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_addr_resize/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_addr_resize/$exit
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_addr_resize/base_resize_req
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_addr_resize/base_resize_ack
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_plus_offset/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_plus_offset/$exit
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_plus_offset/sum_rename_req
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_base_plus_offset/sum_rename_ack
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_sample_start
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_update_start
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_0_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_0_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_0_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_0_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_785/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse43_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse43_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_785/merge_stmt_965_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_785/merge_stmt_965_PhiAck/$entry
      -- CP-element group 79: 	 branch_block_stmt_785/merge_stmt_965_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_785/merge_stmt_965_PhiAck/dummy
      -- 
    if_choice_transition_3530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_959_branch_ack_1, ack => zeropad3D_A_CP_2875_elements(79)); -- 
    cr_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_addr_2_req_1); -- 
    cr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_load_1_req_1); -- 
    rr_3595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_addr_3_req_0); -- 
    cr_3600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_addr_3_req_1); -- 
    rr_3585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_addr_2_req_0); -- 
    cr_3580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_addr_1_req_1); -- 
    cr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_load_0_req_1); -- 
    cr_3652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_load_3_req_1); -- 
    rr_3575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_addr_1_req_0); -- 
    cr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_load_2_req_1); -- 
    rr_3565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_addr_0_req_0); -- 
    cr_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(79), ack => ptr_deref_976_addr_0_req_1); -- 
    -- CP-element group 80:  transition  place  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	77 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	212 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_785/if_stmt_959_else_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_785/if_stmt_959_else_link/else_choice_transition
      -- CP-element group 80: 	 branch_block_stmt_785/lorx_xlhsx_xfalse_ifx_xthen
      -- CP-element group 80: 	 branch_block_stmt_785/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_785/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_959_branch_ack_0, ack => zeropad3D_A_CP_2875_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	92 
    -- CP-element group 81: 	93 
    -- CP-element group 81: 	94 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (11) 
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_3/rr
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_3/$entry
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_2/rr
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_2/$entry
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_1/rr
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_1/$entry
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_0/rr
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/$entry
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_sample_start_
      -- 
    rr_3611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(81), ack => ptr_deref_976_load_0_req_0); -- 
    rr_3616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(81), ack => ptr_deref_976_load_1_req_0); -- 
    rr_3621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(81), ack => ptr_deref_976_load_2_req_0); -- 
    rr_3626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(81), ack => ptr_deref_976_load_3_req_0); -- 
    zeropad3D_A_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(79) & zeropad3D_A_CP_2875_elements(83);
      gj_zeropad3D_A_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: 	86 
    -- CP-element group 82: 	88 
    -- CP-element group 82: 	90 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	102 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_sample_complete
      -- 
    zeropad3D_A_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(84) & zeropad3D_A_CP_2875_elements(86) & zeropad3D_A_CP_2875_elements(88) & zeropad3D_A_CP_2875_elements(90);
      gj_zeropad3D_A_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: 	87 
    -- CP-element group 83: 	89 
    -- CP-element group 83: 	91 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_address_calculated
      -- CP-element group 83: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_update_complete
      -- 
    zeropad3D_A_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(85) & zeropad3D_A_CP_2875_elements(87) & zeropad3D_A_CP_2875_elements(89) & zeropad3D_A_CP_2875_elements(91);
      gj_zeropad3D_A_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	79 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_0_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_0_Sample/ra
      -- 
    ra_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_addr_0_ack_0, ack => zeropad3D_A_CP_2875_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_0_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_0_Update/ca
      -- 
    ca_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_addr_0_ack_1, ack => zeropad3D_A_CP_2875_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	79 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	82 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_1_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_1_Sample/$exit
      -- 
    ra_3576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_addr_1_ack_0, ack => zeropad3D_A_CP_2875_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	79 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	83 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_1_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_1_Update/$exit
      -- 
    ca_3581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_addr_1_ack_1, ack => zeropad3D_A_CP_2875_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	79 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	82 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_2_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_2_Sample/$exit
      -- 
    ra_3586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_addr_2_ack_0, ack => zeropad3D_A_CP_2875_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	79 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	83 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_2_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_2_Update/$exit
      -- 
    ca_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_addr_2_ack_1, ack => zeropad3D_A_CP_2875_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	79 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	82 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_3_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_3_Sample/ra
      -- 
    ra_3596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_addr_3_ack_0, ack => zeropad3D_A_CP_2875_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	79 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	83 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_3_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_word_addrgen_3_Update/ca
      -- 
    ca_3601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_addr_3_ack_1, ack => zeropad3D_A_CP_2875_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	81 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_0/ra
      -- CP-element group 92: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_0/$exit
      -- 
    ra_3612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	81 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	96 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_1/ra
      -- CP-element group 93: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_1/$exit
      -- 
    ra_3617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_load_1_ack_0, ack => zeropad3D_A_CP_2875_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	81 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_2/ra
      -- CP-element group 94: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_2/$exit
      -- 
    ra_3622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_load_2_ack_0, ack => zeropad3D_A_CP_2875_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_3/$exit
      -- CP-element group 95: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/word_3/ra
      -- 
    ra_3627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_load_3_ack_0, ack => zeropad3D_A_CP_2875_elements(95)); -- 
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	93 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/word_access_start/$exit
      -- CP-element group 96: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_sample_completed_
      -- 
    zeropad3D_A_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(92) & zeropad3D_A_CP_2875_elements(93) & zeropad3D_A_CP_2875_elements(94) & zeropad3D_A_CP_2875_elements(95);
      gj_zeropad3D_A_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	79 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_0/ca
      -- CP-element group 97: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_0/$exit
      -- 
    ca_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	79 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	101 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_1/ca
      -- CP-element group 98: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_1/$exit
      -- 
    ca_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_load_1_ack_1, ack => zeropad3D_A_CP_2875_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	79 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_2/ca
      -- CP-element group 99: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_2/$exit
      -- 
    ca_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_load_2_ack_1, ack => zeropad3D_A_CP_2875_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	79 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_3/ca
      -- CP-element group 100: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/word_3/$exit
      -- 
    ca_3653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_976_load_3_ack_1, ack => zeropad3D_A_CP_2875_elements(100)); -- 
    -- CP-element group 101:  join  transition  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: 	97 
    -- CP-element group 101: 	98 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (7) 
      -- CP-element group 101: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/ptr_deref_976_Merge/merge_ack
      -- CP-element group 101: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/ptr_deref_976_Merge/merge_req
      -- CP-element group 101: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/ptr_deref_976_Merge/$exit
      -- CP-element group 101: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/ptr_deref_976_Merge/$entry
      -- CP-element group 101: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/word_access_complete/$exit
      -- CP-element group 101: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/ptr_deref_976_update_completed_
      -- 
    zeropad3D_A_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(99) & zeropad3D_A_CP_2875_elements(100) & zeropad3D_A_CP_2875_elements(97) & zeropad3D_A_CP_2875_elements(98);
      gj_zeropad3D_A_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  branch  join  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: 	82 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (10) 
      -- CP-element group 102: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987__exit__
      -- CP-element group 102: 	 branch_block_stmt_785/if_stmt_988__entry__
      -- CP-element group 102: 	 branch_block_stmt_785/R_cmp49_989_place
      -- CP-element group 102: 	 branch_block_stmt_785/if_stmt_988_else_link/$entry
      -- CP-element group 102: 	 branch_block_stmt_785/if_stmt_988_if_link/$entry
      -- CP-element group 102: 	 branch_block_stmt_785/if_stmt_988_eval_test/branch_req
      -- CP-element group 102: 	 branch_block_stmt_785/if_stmt_988_eval_test/$exit
      -- CP-element group 102: 	 branch_block_stmt_785/if_stmt_988_eval_test/$entry
      -- CP-element group 102: 	 branch_block_stmt_785/if_stmt_988_dead_link/$entry
      -- CP-element group 102: 	 branch_block_stmt_785/assign_stmt_973_to_assign_stmt_987/$exit
      -- 
    branch_req_3666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(102), ack => if_stmt_988_branch_req_0); -- 
    zeropad3D_A_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(101) & zeropad3D_A_CP_2875_elements(82);
      gj_zeropad3D_A_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  place  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	212 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_785/lorx_xlhsx_xfalse43_ifx_xthen
      -- CP-element group 103: 	 branch_block_stmt_785/if_stmt_988_if_link/if_choice_transition
      -- CP-element group 103: 	 branch_block_stmt_785/if_stmt_988_if_link/$exit
      -- CP-element group 103: 	 branch_block_stmt_785/lorx_xlhsx_xfalse43_ifx_xthen_PhiReq/$entry
      -- CP-element group 103: 	 branch_block_stmt_785/lorx_xlhsx_xfalse43_ifx_xthen_PhiReq/$exit
      -- 
    if_choice_transition_3671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_988_branch_ack_1, ack => zeropad3D_A_CP_2875_elements(103)); -- 
    -- CP-element group 104:  fork  transition  place  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	114 
    -- CP-element group 104: 	115 
    -- CP-element group 104: 	117 
    -- CP-element group 104: 	119 
    -- CP-element group 104: 	121 
    -- CP-element group 104: 	122 
    -- CP-element group 104: 	123 
    -- CP-element group 104: 	125 
    -- CP-element group 104: 	127 
    -- CP-element group 104: 	130 
    -- CP-element group 104:  members (46) 
      -- CP-element group 104: 	 branch_block_stmt_785/merge_stmt_1043__exit__
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143__entry__
      -- CP-element group 104: 	 branch_block_stmt_785/lorx_xlhsx_xfalse43_ifx_xelse
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_update_start_
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_complete/req
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_update_start_
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_update_start_
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_785/if_stmt_988_else_link/else_choice_transition
      -- CP-element group 104: 	 branch_block_stmt_785/if_stmt_988_else_link/$exit
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_update_start_
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_update_start_
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_complete/req
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_update_start_
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_785/lorx_xlhsx_xfalse43_ifx_xelse_PhiReq/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/lorx_xlhsx_xfalse43_ifx_xelse_PhiReq/$exit
      -- CP-element group 104: 	 branch_block_stmt_785/merge_stmt_1043_PhiReqMerge
      -- CP-element group 104: 	 branch_block_stmt_785/merge_stmt_1043_PhiAck/$entry
      -- CP-element group 104: 	 branch_block_stmt_785/merge_stmt_1043_PhiAck/$exit
      -- CP-element group 104: 	 branch_block_stmt_785/merge_stmt_1043_PhiAck/dummy
      -- 
    else_choice_transition_3675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_988_branch_ack_0, ack => zeropad3D_A_CP_2875_elements(104)); -- 
    req_3837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => array_obj_ref_1112_index_offset_req_1); -- 
    req_3852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => addr_of_1113_final_reg_req_1); -- 
    cr_3806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => type_cast_1106_inst_req_1); -- 
    rr_3801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => type_cast_1106_inst_req_0); -- 
    cr_3897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => ptr_deref_1117_load_0_req_1); -- 
    rr_3911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => type_cast_1131_inst_req_0); -- 
    cr_3916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => type_cast_1131_inst_req_1); -- 
    req_3947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => array_obj_ref_1137_index_offset_req_1); -- 
    req_3962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => addr_of_1138_final_reg_req_1); -- 
    cr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(104), ack => ptr_deref_1141_store_0_req_1); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	212 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_sample_completed_
      -- 
    ra_3689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1028_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	212 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (16) 
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_resize_1/index_resize_ack
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_resized_1
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_scale_1/$entry
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_scale_1/$exit
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_scale_1/scale_rename_req
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_scale_1/scale_rename_ack
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_scaled_1
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_computed_1
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_resize_1/$entry
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_resize_1/$exit
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_index_resize_1/index_resize_req
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_Sample/req
      -- CP-element group 106: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_Sample/$entry
      -- 
    ca_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1028_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(106)); -- 
    req_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(106), ack => array_obj_ref_1034_index_offset_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	113 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_sample_complete
      -- CP-element group 107: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_Sample/ack
      -- CP-element group 107: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_Sample/$exit
      -- 
    ack_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_offset_ack_0, ack => zeropad3D_A_CP_2875_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	212 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (11) 
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_root_address_calculated
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_offset_calculated
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_request/req
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_request/$entry
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_base_plus_offset/sum_rename_ack
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_base_plus_offset/sum_rename_req
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_base_plus_offset/$exit
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_base_plus_offset/$entry
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_Update/ack
      -- CP-element group 108: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_Update/$exit
      -- 
    ack_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_offset_ack_1, ack => zeropad3D_A_CP_2875_elements(108)); -- 
    req_3734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(108), ack => addr_of_1035_final_reg_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_request/ack
      -- CP-element group 109: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_request/$exit
      -- 
    ack_3735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1035_final_reg_ack_0, ack => zeropad3D_A_CP_2875_elements(109)); -- 
    -- CP-element group 110:  join  fork  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	212 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (28) 
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_addr_resize/base_resize_req
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_plus_offset/$entry
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_addr_resize/base_resize_ack
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_plus_offset/$exit
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_addr_resize/$entry
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_address_resized
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_addr_resize/$exit
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/word_access_start/word_0/$entry
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_plus_offset/sum_rename_req
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_plus_offset/sum_rename_ack
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_word_addrgen/$entry
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/word_access_start/word_0/rr
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_word_addrgen/$exit
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_word_addrgen/root_register_req
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/word_access_start/$entry
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/ptr_deref_1038_Split/split_ack
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/ptr_deref_1038_Split/split_req
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_root_address_calculated
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_word_address_calculated
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/ptr_deref_1038_Split/$exit
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/ptr_deref_1038_Split/$entry
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_base_address_calculated
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_complete/ack
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_word_addrgen/root_register_ack
      -- 
    ack_3740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1035_final_reg_ack_1, ack => zeropad3D_A_CP_2875_elements(110)); -- 
    rr_3778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(110), ack => ptr_deref_1038_store_0_req_0); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/word_access_start/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/word_access_start/word_0/ra
      -- CP-element group 111: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/word_access_start/$exit
      -- CP-element group 111: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Sample/$exit
      -- 
    ra_3779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1038_store_0_ack_0, ack => zeropad3D_A_CP_2875_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	212 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Update/word_access_complete/word_0/ca
      -- CP-element group 112: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Update/word_access_complete/$exit
      -- CP-element group 112: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Update/word_access_complete/word_0/$exit
      -- 
    ca_3790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1038_store_0_ack_1, ack => zeropad3D_A_CP_2875_elements(112)); -- 
    -- CP-element group 113:  join  transition  place  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: 	107 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	213 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041__exit__
      -- CP-element group 113: 	 branch_block_stmt_785/ifx_xthen_ifx_xend
      -- CP-element group 113: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/$exit
      -- CP-element group 113: 	 branch_block_stmt_785/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 113: 	 branch_block_stmt_785/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(112) & zeropad3D_A_CP_2875_elements(107);
      gj_zeropad3D_A_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	104 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_sample_completed_
      -- 
    ra_3802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	104 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (16) 
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_scale_1/$entry
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_scale_1/$exit
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_Sample/req
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_scale_1/scale_rename_req
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_resize_1/index_resize_req
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_scale_1/scale_rename_ack
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_resize_1/index_resize_ack
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_resize_1/$exit
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_resize_1/$entry
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_computed_1
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_scaled_1
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_index_resized_1
      -- CP-element group 115: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1106_Update/$exit
      -- 
    ca_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(115)); -- 
    req_3832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(115), ack => array_obj_ref_1112_index_offset_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	131 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_Sample/ack
      -- CP-element group 116: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_sample_complete
      -- 
    ack_3833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1112_index_offset_ack_0, ack => zeropad3D_A_CP_2875_elements(116)); -- 
    -- CP-element group 117:  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	104 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (11) 
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_root_address_calculated
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_base_plus_offset/sum_rename_ack
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_base_plus_offset/sum_rename_req
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_request/req
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_base_plus_offset/$entry
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_base_plus_offset/$exit
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_request/$entry
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_final_index_sum_regn_Update/ack
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1112_offset_calculated
      -- 
    ack_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1112_index_offset_ack_1, ack => zeropad3D_A_CP_2875_elements(117)); -- 
    req_3847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(117), ack => addr_of_1113_final_reg_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_request/ack
      -- CP-element group 118: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_request/$exit
      -- 
    ack_3848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1113_final_reg_ack_0, ack => zeropad3D_A_CP_2875_elements(118)); -- 
    -- CP-element group 119:  join  fork  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	104 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (24) 
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_complete/$exit
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1113_complete/ack
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Sample/word_access_start/word_0/rr
      -- 
    ack_3853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1113_final_reg_ack_1, ack => zeropad3D_A_CP_2875_elements(119)); -- 
    rr_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(119), ack => ptr_deref_1117_load_0_req_0); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Sample/word_access_start/$exit
      -- CP-element group 120: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Sample/word_access_start/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Sample/word_access_start/word_0/ra
      -- 
    ra_3887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1117_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	104 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	128 
    -- CP-element group 121:  members (9) 
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/word_access_complete/$exit
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/word_access_complete/word_0/$exit
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/word_access_complete/word_0/ca
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/ptr_deref_1117_Merge/$entry
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/ptr_deref_1117_Merge/$exit
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/ptr_deref_1117_Merge/merge_req
      -- CP-element group 121: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1117_Update/ptr_deref_1117_Merge/merge_ack
      -- 
    ca_3898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1117_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	104 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_Sample/ra
      -- 
    ra_3912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1131_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(122)); -- 
    -- CP-element group 123:  transition  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	104 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (16) 
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/type_cast_1131_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_resized_1
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_scaled_1
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_computed_1
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_resize_1/$entry
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_resize_1/$exit
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_resize_1/index_resize_req
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_resize_1/index_resize_ack
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_scale_1/$entry
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_scale_1/$exit
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_scale_1/scale_rename_req
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_index_scale_1/scale_rename_ack
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_Sample/req
      -- 
    ca_3917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1131_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(123)); -- 
    req_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(123), ack => array_obj_ref_1137_index_offset_req_0); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	131 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_sample_complete
      -- CP-element group 124: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_Sample/ack
      -- 
    ack_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1137_index_offset_ack_0, ack => zeropad3D_A_CP_2875_elements(124)); -- 
    -- CP-element group 125:  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	104 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (11) 
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_root_address_calculated
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_offset_calculated
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_final_index_sum_regn_Update/ack
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_base_plus_offset/$entry
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_base_plus_offset/$exit
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_base_plus_offset/sum_rename_req
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/array_obj_ref_1137_base_plus_offset/sum_rename_ack
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_request/$entry
      -- CP-element group 125: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_request/req
      -- 
    ack_3948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1137_index_offset_ack_1, ack => zeropad3D_A_CP_2875_elements(125)); -- 
    req_3957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(125), ack => addr_of_1138_final_reg_req_0); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_request/$exit
      -- CP-element group 126: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_request/ack
      -- 
    ack_3958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1138_final_reg_ack_0, ack => zeropad3D_A_CP_2875_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	104 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (19) 
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_complete/$exit
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/addr_of_1138_complete/ack
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_word_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_root_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_address_resized
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_addr_resize/$entry
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_addr_resize/$exit
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_addr_resize/base_resize_req
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_addr_resize/base_resize_ack
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_plus_offset/$entry
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_plus_offset/$exit
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_plus_offset/sum_rename_req
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_base_plus_offset/sum_rename_ack
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_word_addrgen/$entry
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_word_addrgen/$exit
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_word_addrgen/root_register_req
      -- CP-element group 127: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_word_addrgen/root_register_ack
      -- 
    ack_3963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1138_final_reg_ack_1, ack => zeropad3D_A_CP_2875_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	121 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (9) 
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/ptr_deref_1141_Split/$entry
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/ptr_deref_1141_Split/$exit
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/ptr_deref_1141_Split/split_req
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/ptr_deref_1141_Split/split_ack
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/word_access_start/$entry
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/word_access_start/word_0/$entry
      -- CP-element group 128: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/word_access_start/word_0/rr
      -- 
    rr_4001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(128), ack => ptr_deref_1141_store_0_req_0); -- 
    zeropad3D_A_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(121) & zeropad3D_A_CP_2875_elements(127);
      gj_zeropad3D_A_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/word_access_start/$exit
      -- CP-element group 129: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/word_access_start/word_0/$exit
      -- CP-element group 129: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Sample/word_access_start/word_0/ra
      -- 
    ra_4002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1141_store_0_ack_0, ack => zeropad3D_A_CP_2875_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	104 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (5) 
      -- CP-element group 130: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Update/word_access_complete/$exit
      -- CP-element group 130: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Update/word_access_complete/word_0/$exit
      -- CP-element group 130: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/ptr_deref_1141_Update/word_access_complete/word_0/ca
      -- 
    ca_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1141_store_0_ack_1, ack => zeropad3D_A_CP_2875_elements(130)); -- 
    -- CP-element group 131:  join  transition  place  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	116 
    -- CP-element group 131: 	124 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	213 
    -- CP-element group 131:  members (5) 
      -- CP-element group 131: 	 branch_block_stmt_785/ifx_xelse_ifx_xend
      -- CP-element group 131: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143__exit__
      -- CP-element group 131: 	 branch_block_stmt_785/assign_stmt_1048_to_assign_stmt_1143/$exit
      -- CP-element group 131: 	 branch_block_stmt_785/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 131: 	 branch_block_stmt_785/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(116) & zeropad3D_A_CP_2875_elements(124) & zeropad3D_A_CP_2875_elements(130);
      gj_zeropad3D_A_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  fork  transition  place  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	213 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	214 
    -- CP-element group 132: 	215 
    -- CP-element group 132: 	217 
    -- CP-element group 132: 	218 
    -- CP-element group 132: 	220 
    -- CP-element group 132: 	221 
    -- CP-element group 132:  members (28) 
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116
      -- CP-element group 132: 	 branch_block_stmt_785/if_stmt_1159_if_link/$exit
      -- CP-element group 132: 	 branch_block_stmt_785/if_stmt_1159_if_link/if_choice_transition
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/Update/cr
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/Update/cr
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1159_branch_ack_1, ack => zeropad3D_A_CP_2875_elements(132)); -- 
    rr_4617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(132), ack => type_cast_1220_inst_req_0); -- 
    cr_4622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(132), ack => type_cast_1220_inst_req_1); -- 
    rr_4640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(132), ack => type_cast_1230_inst_req_0); -- 
    cr_4645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(132), ack => type_cast_1230_inst_req_1); -- 
    rr_4663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(132), ack => type_cast_1238_inst_req_0); -- 
    cr_4668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(132), ack => type_cast_1238_inst_req_1); -- 
    -- CP-element group 133:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	213 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133: 	137 
    -- CP-element group 133: 	138 
    -- CP-element group 133: 	139 
    -- CP-element group 133: 	140 
    -- CP-element group 133: 	141 
    -- CP-element group 133: 	142 
    -- CP-element group 133: 	143 
    -- CP-element group 133: 	144 
    -- CP-element group 133: 	150 
    -- CP-element group 133: 	151 
    -- CP-element group 133: 	152 
    -- CP-element group 133: 	153 
    -- CP-element group 133: 	156 
    -- CP-element group 133:  members (55) 
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202__entry__
      -- CP-element group 133: 	 branch_block_stmt_785/merge_stmt_1165__exit__
      -- CP-element group 133: 	 branch_block_stmt_785/ifx_xend_ifx_xthen102
      -- CP-element group 133: 	 branch_block_stmt_785/if_stmt_1159_else_link/$exit
      -- CP-element group 133: 	 branch_block_stmt_785/if_stmt_1159_else_link/else_choice_transition
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_update_start_
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_root_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_address_resized
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_addr_resize/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_addr_resize/$exit
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_addr_resize/base_resize_req
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_addr_resize/base_resize_ack
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_plus_offset/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_plus_offset/$exit
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_plus_offset/sum_rename_req
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_base_plus_offset/sum_rename_ack
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_sample_start
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_update_start
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_0_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_0_Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_0_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_0_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_1_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_1_Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_1_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_1_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_2_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_2_Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_2_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_2_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_3_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_3_Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_3_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_3_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_0/cr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_1/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_1/cr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_2/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_2/cr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_3/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_3/cr
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_update_start_
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_785/ifx_xend_ifx_xthen102_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/ifx_xend_ifx_xthen102_PhiReq/$exit
      -- CP-element group 133: 	 branch_block_stmt_785/merge_stmt_1165_PhiReqMerge
      -- CP-element group 133: 	 branch_block_stmt_785/merge_stmt_1165_PhiAck/$entry
      -- CP-element group 133: 	 branch_block_stmt_785/merge_stmt_1165_PhiAck/$exit
      -- CP-element group 133: 	 branch_block_stmt_785/merge_stmt_1165_PhiAck/dummy
      -- 
    else_choice_transition_4033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1159_branch_ack_0, ack => zeropad3D_A_CP_2875_elements(133)); -- 
    rr_4064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_addr_0_req_0); -- 
    cr_4069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_addr_0_req_1); -- 
    rr_4074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_addr_1_req_0); -- 
    cr_4079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_addr_1_req_1); -- 
    rr_4084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_addr_2_req_0); -- 
    cr_4089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_addr_2_req_1); -- 
    rr_4094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_addr_3_req_0); -- 
    cr_4099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_addr_3_req_1); -- 
    cr_4136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_load_0_req_1); -- 
    cr_4141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_load_1_req_1); -- 
    cr_4146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_load_2_req_1); -- 
    cr_4151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => ptr_deref_1182_load_3_req_1); -- 
    cr_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(133), ack => type_cast_1196_inst_req_1); -- 
    -- CP-element group 134:  join  fork  transition  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: 	136 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	145 
    -- CP-element group 134: 	146 
    -- CP-element group 134: 	147 
    -- CP-element group 134: 	148 
    -- CP-element group 134:  members (11) 
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/$entry
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_0/$entry
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_0/rr
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_1/$entry
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_1/rr
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_2/$entry
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_2/rr
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_3/$entry
      -- CP-element group 134: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_3/rr
      -- 
    rr_4110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(134), ack => ptr_deref_1182_load_0_req_0); -- 
    rr_4115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(134), ack => ptr_deref_1182_load_1_req_0); -- 
    rr_4120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(134), ack => ptr_deref_1182_load_2_req_0); -- 
    rr_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(134), ack => ptr_deref_1182_load_3_req_0); -- 
    zeropad3D_A_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(133) & zeropad3D_A_CP_2875_elements(136);
      gj_zeropad3D_A_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: 	139 
    -- CP-element group 135: 	141 
    -- CP-element group 135: 	143 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	157 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_sample_complete
      -- 
    zeropad3D_A_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(137) & zeropad3D_A_CP_2875_elements(139) & zeropad3D_A_CP_2875_elements(141) & zeropad3D_A_CP_2875_elements(143);
      gj_zeropad3D_A_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: 	140 
    -- CP-element group 136: 	142 
    -- CP-element group 136: 	144 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	134 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_address_calculated
      -- CP-element group 136: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_update_complete
      -- 
    zeropad3D_A_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(138) & zeropad3D_A_CP_2875_elements(140) & zeropad3D_A_CP_2875_elements(142) & zeropad3D_A_CP_2875_elements(144);
      gj_zeropad3D_A_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	133 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	135 
    -- CP-element group 137:  members (2) 
      -- CP-element group 137: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_0_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_0_Sample/ra
      -- 
    ra_4065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_addr_0_ack_0, ack => zeropad3D_A_CP_2875_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	133 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_0_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_0_Update/ca
      -- 
    ca_4070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_addr_0_ack_1, ack => zeropad3D_A_CP_2875_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	133 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	135 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_1_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_1_Sample/ra
      -- 
    ra_4075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_addr_1_ack_0, ack => zeropad3D_A_CP_2875_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	133 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	136 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_1_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_1_Update/ca
      -- 
    ca_4080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_addr_1_ack_1, ack => zeropad3D_A_CP_2875_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	133 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	135 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_2_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_2_Sample/ra
      -- 
    ra_4085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_addr_2_ack_0, ack => zeropad3D_A_CP_2875_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	133 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	136 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_2_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_2_Update/ca
      -- 
    ca_4090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_addr_2_ack_1, ack => zeropad3D_A_CP_2875_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	133 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	135 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_3_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_3_Sample/ra
      -- 
    ra_4095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_addr_3_ack_0, ack => zeropad3D_A_CP_2875_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	133 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	136 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_3_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_word_addrgen_3_Update/ca
      -- 
    ca_4100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_addr_3_ack_1, ack => zeropad3D_A_CP_2875_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	134 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	149 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_0/ra
      -- 
    ra_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	134 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_1/$exit
      -- CP-element group 146: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_1/ra
      -- 
    ra_4116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_load_1_ack_0, ack => zeropad3D_A_CP_2875_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	134 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_2/$exit
      -- CP-element group 147: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_2/ra
      -- 
    ra_4121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_load_2_ack_0, ack => zeropad3D_A_CP_2875_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	134 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_3/$exit
      -- CP-element group 148: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/word_3/ra
      -- 
    ra_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_load_3_ack_0, ack => zeropad3D_A_CP_2875_elements(148)); -- 
    -- CP-element group 149:  join  transition  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	145 
    -- CP-element group 149: 	146 
    -- CP-element group 149: 	147 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Sample/word_access_start/$exit
      -- 
    zeropad3D_A_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(145) & zeropad3D_A_CP_2875_elements(146) & zeropad3D_A_CP_2875_elements(147) & zeropad3D_A_CP_2875_elements(148);
      gj_zeropad3D_A_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	133 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	154 
    -- CP-element group 150:  members (2) 
      -- CP-element group 150: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_0/$exit
      -- CP-element group 150: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_0/ca
      -- 
    ca_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	133 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	154 
    -- CP-element group 151:  members (2) 
      -- CP-element group 151: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_1/$exit
      -- CP-element group 151: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_1/ca
      -- 
    ca_4142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_load_1_ack_1, ack => zeropad3D_A_CP_2875_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	133 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_2/$exit
      -- CP-element group 152: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_2/ca
      -- 
    ca_4147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_load_2_ack_1, ack => zeropad3D_A_CP_2875_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	133 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_3/$exit
      -- CP-element group 153: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/word_3/ca
      -- 
    ca_4152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1182_load_3_ack_1, ack => zeropad3D_A_CP_2875_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	150 
    -- CP-element group 154: 	151 
    -- CP-element group 154: 	152 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (10) 
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/word_access_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/ptr_deref_1182_Merge/$entry
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/ptr_deref_1182_Merge/$exit
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/ptr_deref_1182_Merge/merge_req
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/ptr_deref_1182_Update/ptr_deref_1182_Merge/merge_ack
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_Sample/rr
      -- 
    rr_4165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(154), ack => type_cast_1196_inst_req_0); -- 
    zeropad3D_A_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(150) & zeropad3D_A_CP_2875_elements(151) & zeropad3D_A_CP_2875_elements(152) & zeropad3D_A_CP_2875_elements(153);
      gj_zeropad3D_A_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_Sample/ra
      -- 
    ra_4166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1196_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	133 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/type_cast_1196_Update/ca
      -- 
    ca_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1196_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(156)); -- 
    -- CP-element group 157:  branch  join  transition  place  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	135 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (10) 
      -- CP-element group 157: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202__exit__
      -- CP-element group 157: 	 branch_block_stmt_785/if_stmt_1203__entry__
      -- CP-element group 157: 	 branch_block_stmt_785/assign_stmt_1171_to_assign_stmt_1202/$exit
      -- CP-element group 157: 	 branch_block_stmt_785/if_stmt_1203_dead_link/$entry
      -- CP-element group 157: 	 branch_block_stmt_785/if_stmt_1203_eval_test/$entry
      -- CP-element group 157: 	 branch_block_stmt_785/if_stmt_1203_eval_test/$exit
      -- CP-element group 157: 	 branch_block_stmt_785/if_stmt_1203_eval_test/branch_req
      -- CP-element group 157: 	 branch_block_stmt_785/R_cmp109_1204_place
      -- CP-element group 157: 	 branch_block_stmt_785/if_stmt_1203_if_link/$entry
      -- CP-element group 157: 	 branch_block_stmt_785/if_stmt_1203_else_link/$entry
      -- 
    branch_req_4179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(157), ack => if_stmt_1203_branch_req_0); -- 
    zeropad3D_A_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(135) & zeropad3D_A_CP_2875_elements(156);
      gj_zeropad3D_A_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	232 
    -- CP-element group 158: 	233 
    -- CP-element group 158: 	234 
    -- CP-element group 158: 	235 
    -- CP-element group 158:  members (24) 
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116
      -- CP-element group 158: 	 branch_block_stmt_785/merge_stmt_1209__exit__
      -- CP-element group 158: 	 branch_block_stmt_785/if_stmt_1203_if_link/$exit
      -- CP-element group 158: 	 branch_block_stmt_785/if_stmt_1203_if_link/if_choice_transition
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen102_ifx_xthen111
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen102_ifx_xthen111_PhiReq/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen102_ifx_xthen111_PhiReq/$exit
      -- CP-element group 158: 	 branch_block_stmt_785/merge_stmt_1209_PhiReqMerge
      -- CP-element group 158: 	 branch_block_stmt_785/merge_stmt_1209_PhiAck/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/merge_stmt_1209_PhiAck/$exit
      -- CP-element group 158: 	 branch_block_stmt_785/merge_stmt_1209_PhiAck/dummy
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1212/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1221/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1203_branch_ack_1, ack => zeropad3D_A_CP_2875_elements(158)); -- 
    rr_4762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(158), ack => type_cast_1234_inst_req_0); -- 
    cr_4767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(158), ack => type_cast_1234_inst_req_1); -- 
    -- CP-element group 159:  fork  transition  place  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	224 
    -- CP-element group 159: 	225 
    -- CP-element group 159: 	227 
    -- CP-element group 159: 	228 
    -- CP-element group 159: 	229 
    -- CP-element group 159:  members (22) 
      -- CP-element group 159: 	 branch_block_stmt_785/if_stmt_1203_else_link/$exit
      -- CP-element group 159: 	 branch_block_stmt_785/if_stmt_1203_else_link/else_choice_transition
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/Update/cr
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1221/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1203_branch_ack_0, ack => zeropad3D_A_CP_2875_elements(159)); -- 
    rr_4689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(159), ack => type_cast_1218_inst_req_0); -- 
    cr_4694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(159), ack => type_cast_1218_inst_req_1); -- 
    rr_4720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(159), ack => type_cast_1236_inst_req_0); -- 
    cr_4725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(159), ack => type_cast_1236_inst_req_1); -- 
    -- CP-element group 160:  join  fork  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: 	242 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	171 
    -- CP-element group 160: 	172 
    -- CP-element group 160: 	173 
    -- CP-element group 160: 	174 
    -- CP-element group 160:  members (11) 
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/$entry
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_0/$entry
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_0/rr
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_1/$entry
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_1/rr
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_2/$entry
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_2/rr
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_3/$entry
      -- CP-element group 160: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_3/rr
      -- 
    rr_4265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(160), ack => ptr_deref_1250_load_0_req_0); -- 
    rr_4270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(160), ack => ptr_deref_1250_load_1_req_0); -- 
    rr_4275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(160), ack => ptr_deref_1250_load_2_req_0); -- 
    rr_4280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(160), ack => ptr_deref_1250_load_3_req_0); -- 
    zeropad3D_A_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(162) & zeropad3D_A_CP_2875_elements(242);
      gj_zeropad3D_A_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	165 
    -- CP-element group 161: 	167 
    -- CP-element group 161: 	169 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	181 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_sample_complete
      -- 
    zeropad3D_A_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(163) & zeropad3D_A_CP_2875_elements(165) & zeropad3D_A_CP_2875_elements(167) & zeropad3D_A_CP_2875_elements(169);
      gj_zeropad3D_A_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  join  transition  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: 	166 
    -- CP-element group 162: 	168 
    -- CP-element group 162: 	170 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_address_calculated
      -- CP-element group 162: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_update_complete
      -- 
    zeropad3D_A_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(164) & zeropad3D_A_CP_2875_elements(166) & zeropad3D_A_CP_2875_elements(168) & zeropad3D_A_CP_2875_elements(170);
      gj_zeropad3D_A_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	242 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_0_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_0_Sample/ra
      -- 
    ra_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_addr_0_ack_0, ack => zeropad3D_A_CP_2875_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	242 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_0_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_0_Update/ca
      -- 
    ca_4225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_addr_0_ack_1, ack => zeropad3D_A_CP_2875_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	242 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	161 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_1_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_1_Sample/ra
      -- 
    ra_4230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_addr_1_ack_0, ack => zeropad3D_A_CP_2875_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	242 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	162 
    -- CP-element group 166:  members (2) 
      -- CP-element group 166: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_1_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_1_Update/ca
      -- 
    ca_4235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_addr_1_ack_1, ack => zeropad3D_A_CP_2875_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	242 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	161 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_2_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_2_Sample/ra
      -- 
    ra_4240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_addr_2_ack_0, ack => zeropad3D_A_CP_2875_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	242 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	162 
    -- CP-element group 168:  members (2) 
      -- CP-element group 168: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_2_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_2_Update/ca
      -- 
    ca_4245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_addr_2_ack_1, ack => zeropad3D_A_CP_2875_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	242 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	161 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_3_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_3_Sample/ra
      -- 
    ra_4250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_addr_3_ack_0, ack => zeropad3D_A_CP_2875_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	242 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	162 
    -- CP-element group 170:  members (2) 
      -- CP-element group 170: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_3_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_3_Update/ca
      -- 
    ca_4255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_addr_3_ack_1, ack => zeropad3D_A_CP_2875_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	160 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	175 
    -- CP-element group 171:  members (2) 
      -- CP-element group 171: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_0/$exit
      -- CP-element group 171: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_0/ra
      -- 
    ra_4266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_0_ack_0, ack => zeropad3D_A_CP_2875_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	160 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	175 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_1/$exit
      -- CP-element group 172: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_1/ra
      -- 
    ra_4271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_1_ack_0, ack => zeropad3D_A_CP_2875_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	160 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (2) 
      -- CP-element group 173: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_2/$exit
      -- CP-element group 173: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_2/ra
      -- 
    ra_4276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_2_ack_0, ack => zeropad3D_A_CP_2875_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	160 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (2) 
      -- CP-element group 174: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_3/$exit
      -- CP-element group 174: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/word_3/ra
      -- 
    ra_4281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_3_ack_0, ack => zeropad3D_A_CP_2875_elements(174)); -- 
    -- CP-element group 175:  join  transition  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	171 
    -- CP-element group 175: 	172 
    -- CP-element group 175: 	173 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Sample/word_access_start/$exit
      -- 
    zeropad3D_A_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(171) & zeropad3D_A_CP_2875_elements(172) & zeropad3D_A_CP_2875_elements(173) & zeropad3D_A_CP_2875_elements(174);
      gj_zeropad3D_A_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	242 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	180 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_0/$exit
      -- CP-element group 176: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_0/ca
      -- 
    ca_4292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_0_ack_1, ack => zeropad3D_A_CP_2875_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	242 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	180 
    -- CP-element group 177:  members (2) 
      -- CP-element group 177: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_1/$exit
      -- CP-element group 177: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_1/ca
      -- 
    ca_4297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_1_ack_1, ack => zeropad3D_A_CP_2875_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	242 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_2/$exit
      -- CP-element group 178: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_2/ca
      -- 
    ca_4302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_2_ack_1, ack => zeropad3D_A_CP_2875_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	242 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_3/$exit
      -- CP-element group 179: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_3/ca
      -- 
    ca_4307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1250_load_3_ack_1, ack => zeropad3D_A_CP_2875_elements(179)); -- 
    -- CP-element group 180:  join  transition  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	176 
    -- CP-element group 180: 	177 
    -- CP-element group 180: 	178 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (7) 
      -- CP-element group 180: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/$exit
      -- CP-element group 180: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/ptr_deref_1250_Merge/$entry
      -- CP-element group 180: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/ptr_deref_1250_Merge/$exit
      -- CP-element group 180: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/ptr_deref_1250_Merge/merge_req
      -- CP-element group 180: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/ptr_deref_1250_Merge/merge_ack
      -- 
    zeropad3D_A_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(176) & zeropad3D_A_CP_2875_elements(177) & zeropad3D_A_CP_2875_elements(178) & zeropad3D_A_CP_2875_elements(179);
      gj_zeropad3D_A_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  branch  join  transition  place  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: 	161 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (10) 
      -- CP-element group 181: 	 branch_block_stmt_785/if_stmt_1262__entry__
      -- CP-element group 181: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261__exit__
      -- CP-element group 181: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/$exit
      -- CP-element group 181: 	 branch_block_stmt_785/if_stmt_1262_dead_link/$entry
      -- CP-element group 181: 	 branch_block_stmt_785/if_stmt_1262_eval_test/$entry
      -- CP-element group 181: 	 branch_block_stmt_785/if_stmt_1262_eval_test/$exit
      -- CP-element group 181: 	 branch_block_stmt_785/if_stmt_1262_eval_test/branch_req
      -- CP-element group 181: 	 branch_block_stmt_785/R_cmp_1263_place
      -- CP-element group 181: 	 branch_block_stmt_785/if_stmt_1262_if_link/$entry
      -- CP-element group 181: 	 branch_block_stmt_785/if_stmt_1262_else_link/$entry
      -- 
    branch_req_4320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(181), ack => if_stmt_1262_branch_req_0); -- 
    zeropad3D_A_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(180) & zeropad3D_A_CP_2875_elements(161);
      gj_zeropad3D_A_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  place  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	193 
    -- CP-element group 182: 	194 
    -- CP-element group 182: 	196 
    -- CP-element group 182: 	197 
    -- CP-element group 182: 	199 
    -- CP-element group 182: 	200 
    -- CP-element group 182: 	202 
    -- CP-element group 182: 	203 
    -- CP-element group 182:  members (36) 
      -- CP-element group 182: 	 branch_block_stmt_785/if_stmt_1262_if_link/$exit
      -- CP-element group 182: 	 branch_block_stmt_785/if_stmt_1262_if_link/if_choice_transition
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/Update/cr
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/Update/cr
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/Update/cr
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1262_branch_ack_1, ack => zeropad3D_A_CP_2875_elements(182)); -- 
    rr_4429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(182), ack => type_cast_899_inst_req_0); -- 
    cr_4434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(182), ack => type_cast_899_inst_req_1); -- 
    rr_4452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(182), ack => type_cast_906_inst_req_0); -- 
    cr_4457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(182), ack => type_cast_906_inst_req_1); -- 
    rr_4475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(182), ack => type_cast_913_inst_req_0); -- 
    cr_4480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(182), ack => type_cast_913_inst_req_1); -- 
    rr_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(182), ack => type_cast_920_inst_req_0); -- 
    cr_4503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(182), ack => type_cast_920_inst_req_1); -- 
    -- CP-element group 183:  merge  transition  place  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	243 
    -- CP-element group 183:  members (13) 
      -- CP-element group 183: 	 branch_block_stmt_785/whilex_xendx_xloopexit_whilex_xend
      -- CP-element group 183: 	 branch_block_stmt_785/merge_stmt_1268__exit__
      -- CP-element group 183: 	 branch_block_stmt_785/if_stmt_1262_else_link/$exit
      -- CP-element group 183: 	 branch_block_stmt_785/if_stmt_1262_else_link/else_choice_transition
      -- CP-element group 183: 	 branch_block_stmt_785/ifx_xend116_whilex_xendx_xloopexit
      -- CP-element group 183: 	 branch_block_stmt_785/whilex_xendx_xloopexit_whilex_xend_PhiReq/$exit
      -- CP-element group 183: 	 branch_block_stmt_785/whilex_xendx_xloopexit_whilex_xend_PhiReq/$entry
      -- CP-element group 183: 	 branch_block_stmt_785/merge_stmt_1268_PhiAck/dummy
      -- CP-element group 183: 	 branch_block_stmt_785/ifx_xend116_whilex_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 183: 	 branch_block_stmt_785/ifx_xend116_whilex_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 183: 	 branch_block_stmt_785/merge_stmt_1268_PhiReqMerge
      -- CP-element group 183: 	 branch_block_stmt_785/merge_stmt_1268_PhiAck/$entry
      -- CP-element group 183: 	 branch_block_stmt_785/merge_stmt_1268_PhiAck/$exit
      -- 
    else_choice_transition_4329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1262_branch_ack_0, ack => zeropad3D_A_CP_2875_elements(183)); -- 
    -- CP-element group 184:  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	243 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (6) 
      -- CP-element group 184: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_update_start_
      -- CP-element group 184: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_Sample/ack
      -- CP-element group 184: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_Update/req
      -- 
    ack_4343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1272_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(184)); -- 
    req_4347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(184), ack => WPIPE_Block0_complete_1272_inst_req_1); -- 
    -- CP-element group 185:  transition  place  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (16) 
      -- CP-element group 185: 	 branch_block_stmt_785/branch_block_stmt_785__exit__
      -- CP-element group 185: 	 branch_block_stmt_785/return__
      -- CP-element group 185: 	 branch_block_stmt_785/assign_stmt_1274__exit__
      -- CP-element group 185: 	 branch_block_stmt_785/$exit
      -- CP-element group 185: 	 branch_block_stmt_785/merge_stmt_1276__exit__
      -- CP-element group 185: 	 $exit
      -- CP-element group 185: 	 branch_block_stmt_785/merge_stmt_1276_PhiAck/dummy
      -- CP-element group 185: 	 branch_block_stmt_785/merge_stmt_1276_PhiReqMerge
      -- CP-element group 185: 	 branch_block_stmt_785/return___PhiReq/$exit
      -- CP-element group 185: 	 branch_block_stmt_785/merge_stmt_1276_PhiAck/$entry
      -- CP-element group 185: 	 branch_block_stmt_785/merge_stmt_1276_PhiAck/$exit
      -- CP-element group 185: 	 branch_block_stmt_785/return___PhiReq/$entry
      -- CP-element group 185: 	 branch_block_stmt_785/assign_stmt_1274/$exit
      -- CP-element group 185: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_Update/ack
      -- 
    ack_4348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1272_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	76 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (2) 
      -- CP-element group 186: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/Sample/ra
      -- 
    ra_4380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(186)); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	76 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (2) 
      -- CP-element group 187: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/Update/ca
      -- 
    ca_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	192 
    -- CP-element group 188:  members (5) 
      -- CP-element group 188: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/$exit
      -- CP-element group 188: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/$exit
      -- CP-element group 188: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/$exit
      -- CP-element group 188: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897/SplitProtocol/$exit
      -- CP-element group 188: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_req
      -- 
    phi_stmt_894_req_4386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_894_req_4386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(188), ack => phi_stmt_894_req_0); -- 
    zeropad3D_A_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(186) & zeropad3D_A_CP_2875_elements(187);
      gj_zeropad3D_A_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  transition  output  delay-element  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	76 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	192 
    -- CP-element group 189:  members (4) 
      -- CP-element group 189: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_900/$exit
      -- CP-element group 189: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/$exit
      -- CP-element group 189: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_904_konst_delay_trans
      -- CP-element group 189: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_req
      -- 
    phi_stmt_900_req_4394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_900_req_4394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(189), ack => phi_stmt_900_req_0); -- 
    -- Element group zeropad3D_A_CP_2875_elements(189) is a control-delay.
    cp_element_189_delay: control_delay_element  generic map(name => " 189_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2875_elements(76), ack => zeropad3D_A_CP_2875_elements(189), clk => clk, reset =>reset);
    -- CP-element group 190:  transition  output  delay-element  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	76 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (4) 
      -- CP-element group 190: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_907/$exit
      -- CP-element group 190: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/$exit
      -- CP-element group 190: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_911_konst_delay_trans
      -- CP-element group 190: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_req
      -- 
    phi_stmt_907_req_4402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_907_req_4402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(190), ack => phi_stmt_907_req_0); -- 
    -- Element group zeropad3D_A_CP_2875_elements(190) is a control-delay.
    cp_element_190_delay: control_delay_element  generic map(name => " 190_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2875_elements(76), ack => zeropad3D_A_CP_2875_elements(190), clk => clk, reset =>reset);
    -- CP-element group 191:  transition  output  delay-element  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	76 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (4) 
      -- CP-element group 191: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_914/$exit
      -- CP-element group 191: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/$exit
      -- CP-element group 191: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_918_konst_delay_trans
      -- CP-element group 191: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_req
      -- 
    phi_stmt_914_req_4410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_914_req_4410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(191), ack => phi_stmt_914_req_0); -- 
    -- Element group zeropad3D_A_CP_2875_elements(191) is a control-delay.
    cp_element_191_delay: control_delay_element  generic map(name => " 191_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2875_elements(76), ack => zeropad3D_A_CP_2875_elements(191), clk => clk, reset =>reset);
    -- CP-element group 192:  join  transition  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: 	191 
    -- CP-element group 192: 	189 
    -- CP-element group 192: 	188 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	206 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_785/bbx_xnph_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(190) & zeropad3D_A_CP_2875_elements(191) & zeropad3D_A_CP_2875_elements(189) & zeropad3D_A_CP_2875_elements(188);
      gj_zeropad3D_A_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	182 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (2) 
      -- CP-element group 193: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/Sample/ra
      -- 
    ra_4430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_899_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	182 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (2) 
      -- CP-element group 194: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/Update/ca
      -- 
    ca_4435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_899_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	205 
    -- CP-element group 195:  members (5) 
      -- CP-element group 195: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/$exit
      -- CP-element group 195: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/$exit
      -- CP-element group 195: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/$exit
      -- CP-element group 195: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_899/SplitProtocol/$exit
      -- CP-element group 195: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_894/phi_stmt_894_req
      -- 
    phi_stmt_894_req_4436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_894_req_4436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(195), ack => phi_stmt_894_req_1); -- 
    zeropad3D_A_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(193) & zeropad3D_A_CP_2875_elements(194);
      gj_zeropad3D_A_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	182 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (2) 
      -- CP-element group 196: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/Sample/ra
      -- 
    ra_4453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_906_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	182 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/Update/ca
      -- 
    ca_4458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_906_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	205 
    -- CP-element group 198:  members (5) 
      -- CP-element group 198: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/$exit
      -- CP-element group 198: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/$exit
      -- CP-element group 198: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/$exit
      -- CP-element group 198: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906/SplitProtocol/$exit
      -- CP-element group 198: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_900/phi_stmt_900_req
      -- 
    phi_stmt_900_req_4459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_900_req_4459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(198), ack => phi_stmt_900_req_1); -- 
    zeropad3D_A_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(196) & zeropad3D_A_CP_2875_elements(197);
      gj_zeropad3D_A_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	182 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/Sample/ra
      -- 
    ra_4476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_913_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	182 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (2) 
      -- CP-element group 200: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/Update/ca
      -- 
    ca_4481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_913_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(200)); -- 
    -- CP-element group 201:  join  transition  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	205 
    -- CP-element group 201:  members (5) 
      -- CP-element group 201: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/$exit
      -- CP-element group 201: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/$exit
      -- CP-element group 201: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/$exit
      -- CP-element group 201: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_sources/type_cast_913/SplitProtocol/$exit
      -- CP-element group 201: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_907/phi_stmt_907_req
      -- 
    phi_stmt_907_req_4482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_907_req_4482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(201), ack => phi_stmt_907_req_1); -- 
    zeropad3D_A_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(199) & zeropad3D_A_CP_2875_elements(200);
      gj_zeropad3D_A_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	182 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/Sample/ra
      -- 
    ra_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_920_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(202)); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	182 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (2) 
      -- CP-element group 203: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/Update/ca
      -- 
    ca_4504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_920_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/$exit
      -- CP-element group 204: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/$exit
      -- CP-element group 204: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/$exit
      -- CP-element group 204: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_sources/type_cast_920/SplitProtocol/$exit
      -- CP-element group 204: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/phi_stmt_914/phi_stmt_914_req
      -- 
    phi_stmt_914_req_4505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_914_req_4505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(204), ack => phi_stmt_914_req_1); -- 
    zeropad3D_A_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(202) & zeropad3D_A_CP_2875_elements(203);
      gj_zeropad3D_A_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  join  transition  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	195 
    -- CP-element group 205: 	198 
    -- CP-element group 205: 	201 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_785/ifx_xend116_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(195) & zeropad3D_A_CP_2875_elements(198) & zeropad3D_A_CP_2875_elements(201) & zeropad3D_A_CP_2875_elements(204);
      gj_zeropad3D_A_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  merge  fork  transition  place  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	192 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: 	208 
    -- CP-element group 206: 	209 
    -- CP-element group 206: 	210 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_785/merge_stmt_893_PhiReqMerge
      -- CP-element group 206: 	 branch_block_stmt_785/merge_stmt_893_PhiAck/$entry
      -- 
    zeropad3D_A_CP_2875_elements(206) <= OrReduce(zeropad3D_A_CP_2875_elements(192) & zeropad3D_A_CP_2875_elements(205));
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	211 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_785/merge_stmt_893_PhiAck/phi_stmt_894_ack
      -- 
    phi_stmt_894_ack_4510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_894_ack_0, ack => zeropad3D_A_CP_2875_elements(207)); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	211 
    -- CP-element group 208:  members (1) 
      -- CP-element group 208: 	 branch_block_stmt_785/merge_stmt_893_PhiAck/phi_stmt_900_ack
      -- 
    phi_stmt_900_ack_4511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_900_ack_0, ack => zeropad3D_A_CP_2875_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	206 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_785/merge_stmt_893_PhiAck/phi_stmt_907_ack
      -- 
    phi_stmt_907_ack_4512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_907_ack_0, ack => zeropad3D_A_CP_2875_elements(209)); -- 
    -- CP-element group 210:  transition  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	206 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_785/merge_stmt_893_PhiAck/phi_stmt_914_ack
      -- 
    phi_stmt_914_ack_4513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_914_ack_0, ack => zeropad3D_A_CP_2875_elements(210)); -- 
    -- CP-element group 211:  branch  join  transition  place  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	207 
    -- CP-element group 211: 	208 
    -- CP-element group 211: 	209 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	77 
    -- CP-element group 211: 	78 
    -- CP-element group 211:  members (14) 
      -- CP-element group 211: 	 branch_block_stmt_785/merge_stmt_893__exit__
      -- CP-element group 211: 	 branch_block_stmt_785/assign_stmt_929__entry__
      -- CP-element group 211: 	 branch_block_stmt_785/assign_stmt_929__exit__
      -- CP-element group 211: 	 branch_block_stmt_785/if_stmt_930__entry__
      -- CP-element group 211: 	 branch_block_stmt_785/assign_stmt_929/$entry
      -- CP-element group 211: 	 branch_block_stmt_785/assign_stmt_929/$exit
      -- CP-element group 211: 	 branch_block_stmt_785/if_stmt_930_dead_link/$entry
      -- CP-element group 211: 	 branch_block_stmt_785/if_stmt_930_eval_test/$entry
      -- CP-element group 211: 	 branch_block_stmt_785/if_stmt_930_eval_test/$exit
      -- CP-element group 211: 	 branch_block_stmt_785/if_stmt_930_eval_test/branch_req
      -- CP-element group 211: 	 branch_block_stmt_785/R_cmp28_931_place
      -- CP-element group 211: 	 branch_block_stmt_785/if_stmt_930_if_link/$entry
      -- CP-element group 211: 	 branch_block_stmt_785/if_stmt_930_else_link/$entry
      -- CP-element group 211: 	 branch_block_stmt_785/merge_stmt_893_PhiAck/$exit
      -- 
    branch_req_3503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(211), ack => if_stmt_930_branch_req_0); -- 
    zeropad3D_A_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(207) & zeropad3D_A_CP_2875_elements(208) & zeropad3D_A_CP_2875_elements(209) & zeropad3D_A_CP_2875_elements(210);
      gj_zeropad3D_A_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  merge  fork  transition  place  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	103 
    -- CP-element group 212: 	78 
    -- CP-element group 212: 	80 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	110 
    -- CP-element group 212: 	112 
    -- CP-element group 212: 	105 
    -- CP-element group 212: 	108 
    -- CP-element group 212: 	106 
    -- CP-element group 212:  members (24) 
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041__entry__
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_update_start_
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_update_start
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Update/word_access_complete/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/merge_stmt_994__exit__
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_Update/cr
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_update_start_
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_complete/req
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/addr_of_1035_complete/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_update_start_
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Update/word_access_complete/word_0/cr
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/type_cast_1028_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_Update/req
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/array_obj_ref_1034_final_index_sum_regn_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/assign_stmt_999_to_assign_stmt_1041/ptr_deref_1038_Update/word_access_complete/word_0/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/merge_stmt_994_PhiReqMerge
      -- CP-element group 212: 	 branch_block_stmt_785/merge_stmt_994_PhiAck/$entry
      -- CP-element group 212: 	 branch_block_stmt_785/merge_stmt_994_PhiAck/$exit
      -- CP-element group 212: 	 branch_block_stmt_785/merge_stmt_994_PhiAck/dummy
      -- 
    cr_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(212), ack => type_cast_1028_inst_req_1); -- 
    rr_3688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(212), ack => type_cast_1028_inst_req_0); -- 
    req_3739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(212), ack => addr_of_1035_final_reg_req_1); -- 
    cr_3789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(212), ack => ptr_deref_1038_store_0_req_1); -- 
    req_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(212), ack => array_obj_ref_1034_index_offset_req_1); -- 
    zeropad3D_A_CP_2875_elements(212) <= OrReduce(zeropad3D_A_CP_2875_elements(103) & zeropad3D_A_CP_2875_elements(78) & zeropad3D_A_CP_2875_elements(80));
    -- CP-element group 213:  merge  branch  transition  place  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	113 
    -- CP-element group 213: 	131 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	132 
    -- CP-element group 213: 	133 
    -- CP-element group 213:  members (17) 
      -- CP-element group 213: 	 branch_block_stmt_785/merge_stmt_1145__exit__
      -- CP-element group 213: 	 branch_block_stmt_785/R_cmp100_1160_place
      -- CP-element group 213: 	 branch_block_stmt_785/assign_stmt_1151_to_assign_stmt_1158__entry__
      -- CP-element group 213: 	 branch_block_stmt_785/assign_stmt_1151_to_assign_stmt_1158__exit__
      -- CP-element group 213: 	 branch_block_stmt_785/if_stmt_1159__entry__
      -- CP-element group 213: 	 branch_block_stmt_785/assign_stmt_1151_to_assign_stmt_1158/$entry
      -- CP-element group 213: 	 branch_block_stmt_785/assign_stmt_1151_to_assign_stmt_1158/$exit
      -- CP-element group 213: 	 branch_block_stmt_785/if_stmt_1159_dead_link/$entry
      -- CP-element group 213: 	 branch_block_stmt_785/if_stmt_1159_eval_test/$entry
      -- CP-element group 213: 	 branch_block_stmt_785/if_stmt_1159_eval_test/$exit
      -- CP-element group 213: 	 branch_block_stmt_785/if_stmt_1159_eval_test/branch_req
      -- CP-element group 213: 	 branch_block_stmt_785/if_stmt_1159_if_link/$entry
      -- CP-element group 213: 	 branch_block_stmt_785/if_stmt_1159_else_link/$entry
      -- CP-element group 213: 	 branch_block_stmt_785/merge_stmt_1145_PhiReqMerge
      -- CP-element group 213: 	 branch_block_stmt_785/merge_stmt_1145_PhiAck/$entry
      -- CP-element group 213: 	 branch_block_stmt_785/merge_stmt_1145_PhiAck/$exit
      -- CP-element group 213: 	 branch_block_stmt_785/merge_stmt_1145_PhiAck/dummy
      -- 
    branch_req_4024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(213), ack => if_stmt_1159_branch_req_0); -- 
    zeropad3D_A_CP_2875_elements(213) <= OrReduce(zeropad3D_A_CP_2875_elements(113) & zeropad3D_A_CP_2875_elements(131));
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	132 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (2) 
      -- CP-element group 214: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/Sample/ra
      -- 
    ra_4618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	132 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (2) 
      -- CP-element group 215: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/Update/ca
      -- 
    ca_4623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	223 
    -- CP-element group 216:  members (5) 
      -- CP-element group 216: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/$exit
      -- CP-element group 216: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/$exit
      -- CP-element group 216: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/$exit
      -- CP-element group 216: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1220/SplitProtocol/$exit
      -- CP-element group 216: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_req
      -- 
    phi_stmt_1212_req_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1212_req_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(216), ack => phi_stmt_1212_req_2); -- 
    zeropad3D_A_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(214) & zeropad3D_A_CP_2875_elements(215);
      gj_zeropad3D_A_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	132 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/Sample/ra
      -- 
    ra_4641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	132 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/Update/ca
      -- 
    ca_4646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	223 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/$exit
      -- CP-element group 219: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/$exit
      -- CP-element group 219: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/$exit
      -- CP-element group 219: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1230/SplitProtocol/$exit
      -- CP-element group 219: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_req
      -- 
    phi_stmt_1221_req_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1221_req_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(219), ack => phi_stmt_1221_req_2); -- 
    zeropad3D_A_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(217) & zeropad3D_A_CP_2875_elements(218);
      gj_zeropad3D_A_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	132 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/Sample/ra
      -- 
    ra_4664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	132 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (2) 
      -- CP-element group 221: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/Update/ca
      -- 
    ca_4669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (5) 
      -- CP-element group 222: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/$exit
      -- CP-element group 222: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/$exit
      -- CP-element group 222: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/$exit
      -- CP-element group 222: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1238/SplitProtocol/$exit
      -- CP-element group 222: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_req
      -- 
    phi_stmt_1231_req_4670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1231_req_4670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(222), ack => phi_stmt_1231_req_2); -- 
    zeropad3D_A_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(220) & zeropad3D_A_CP_2875_elements(221);
      gj_zeropad3D_A_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	216 
    -- CP-element group 223: 	219 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	238 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_785/ifx_xend_ifx_xend116_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(216) & zeropad3D_A_CP_2875_elements(219) & zeropad3D_A_CP_2875_elements(222);
      gj_zeropad3D_A_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	159 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	226 
    -- CP-element group 224:  members (2) 
      -- CP-element group 224: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/Sample/ra
      -- 
    ra_4690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	159 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/Update/ca
      -- 
    ca_4695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	231 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/$exit
      -- CP-element group 226: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/$exit
      -- CP-element group 226: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/$exit
      -- CP-element group 226: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1218/SplitProtocol/$exit
      -- CP-element group 226: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_req
      -- 
    phi_stmt_1212_req_4696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1212_req_4696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(226), ack => phi_stmt_1212_req_1); -- 
    zeropad3D_A_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(224) & zeropad3D_A_CP_2875_elements(225);
      gj_zeropad3D_A_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  transition  output  delay-element  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	159 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	231 
    -- CP-element group 227:  members (4) 
      -- CP-element group 227: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1221/$exit
      -- CP-element group 227: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/$exit
      -- CP-element group 227: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1228_konst_delay_trans
      -- CP-element group 227: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_req
      -- 
    phi_stmt_1221_req_4704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1221_req_4704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(227), ack => phi_stmt_1221_req_1); -- 
    -- Element group zeropad3D_A_CP_2875_elements(227) is a control-delay.
    cp_element_227_delay: control_delay_element  generic map(name => " 227_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2875_elements(159), ack => zeropad3D_A_CP_2875_elements(227), clk => clk, reset =>reset);
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	159 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/Sample/ra
      -- 
    ra_4721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1236_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	159 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (2) 
      -- CP-element group 229: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/Update/ca
      -- 
    ca_4726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1236_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/$exit
      -- CP-element group 230: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/$exit
      -- CP-element group 230: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/$exit
      -- CP-element group 230: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1236/SplitProtocol/$exit
      -- CP-element group 230: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_req
      -- 
    phi_stmt_1231_req_4727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1231_req_4727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(230), ack => phi_stmt_1231_req_1); -- 
    zeropad3D_A_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(228) & zeropad3D_A_CP_2875_elements(229);
      gj_zeropad3D_A_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	226 
    -- CP-element group 231: 	227 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	238 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 branch_block_stmt_785/ifx_xthen102_ifx_xend116_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(226) & zeropad3D_A_CP_2875_elements(227) & zeropad3D_A_CP_2875_elements(230);
      gj_zeropad3D_A_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  transition  output  delay-element  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	158 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	237 
    -- CP-element group 232:  members (4) 
      -- CP-element group 232: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1212/$exit
      -- CP-element group 232: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/$exit
      -- CP-element group 232: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_sources/type_cast_1216_konst_delay_trans
      -- CP-element group 232: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1212/phi_stmt_1212_req
      -- 
    phi_stmt_1212_req_4738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1212_req_4738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(232), ack => phi_stmt_1212_req_0); -- 
    -- Element group zeropad3D_A_CP_2875_elements(232) is a control-delay.
    cp_element_232_delay: control_delay_element  generic map(name => " 232_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2875_elements(158), ack => zeropad3D_A_CP_2875_elements(232), clk => clk, reset =>reset);
    -- CP-element group 233:  transition  output  delay-element  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	158 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	237 
    -- CP-element group 233:  members (4) 
      -- CP-element group 233: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1221/$exit
      -- CP-element group 233: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/$exit
      -- CP-element group 233: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_sources/type_cast_1225_konst_delay_trans
      -- CP-element group 233: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1221/phi_stmt_1221_req
      -- 
    phi_stmt_1221_req_4746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1221_req_4746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(233), ack => phi_stmt_1221_req_0); -- 
    -- Element group zeropad3D_A_CP_2875_elements(233) is a control-delay.
    cp_element_233_delay: control_delay_element  generic map(name => " 233_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_2875_elements(158), ack => zeropad3D_A_CP_2875_elements(233), clk => clk, reset =>reset);
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	158 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/Sample/ra
      -- 
    ra_4763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_0, ack => zeropad3D_A_CP_2875_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	158 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/Update/ca
      -- 
    ca_4768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_1, ack => zeropad3D_A_CP_2875_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (5) 
      -- CP-element group 236: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/$exit
      -- CP-element group 236: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/$exit
      -- CP-element group 236: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/$exit
      -- CP-element group 236: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_sources/type_cast_1234/SplitProtocol/$exit
      -- CP-element group 236: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/phi_stmt_1231/phi_stmt_1231_req
      -- 
    phi_stmt_1231_req_4769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1231_req_4769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(236), ack => phi_stmt_1231_req_0); -- 
    zeropad3D_A_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(234) & zeropad3D_A_CP_2875_elements(235);
      gj_zeropad3D_A_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	232 
    -- CP-element group 237: 	233 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (1) 
      -- CP-element group 237: 	 branch_block_stmt_785/ifx_xthen111_ifx_xend116_PhiReq/$exit
      -- 
    zeropad3D_A_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(232) & zeropad3D_A_CP_2875_elements(233) & zeropad3D_A_CP_2875_elements(236);
      gj_zeropad3D_A_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  merge  fork  transition  place  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	223 
    -- CP-element group 238: 	231 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: 	240 
    -- CP-element group 238: 	241 
    -- CP-element group 238:  members (2) 
      -- CP-element group 238: 	 branch_block_stmt_785/merge_stmt_1211_PhiReqMerge
      -- CP-element group 238: 	 branch_block_stmt_785/merge_stmt_1211_PhiAck/$entry
      -- 
    zeropad3D_A_CP_2875_elements(238) <= OrReduce(zeropad3D_A_CP_2875_elements(223) & zeropad3D_A_CP_2875_elements(231) & zeropad3D_A_CP_2875_elements(237));
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	242 
    -- CP-element group 239:  members (1) 
      -- CP-element group 239: 	 branch_block_stmt_785/merge_stmt_1211_PhiAck/phi_stmt_1212_ack
      -- 
    phi_stmt_1212_ack_4774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1212_ack_0, ack => zeropad3D_A_CP_2875_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (1) 
      -- CP-element group 240: 	 branch_block_stmt_785/merge_stmt_1211_PhiAck/phi_stmt_1221_ack
      -- 
    phi_stmt_1221_ack_4775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1221_ack_0, ack => zeropad3D_A_CP_2875_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	238 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (1) 
      -- CP-element group 241: 	 branch_block_stmt_785/merge_stmt_1211_PhiAck/phi_stmt_1231_ack
      -- 
    phi_stmt_1231_ack_4776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1231_ack_0, ack => zeropad3D_A_CP_2875_elements(241)); -- 
    -- CP-element group 242:  join  fork  transition  place  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	239 
    -- CP-element group 242: 	240 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	160 
    -- CP-element group 242: 	163 
    -- CP-element group 242: 	164 
    -- CP-element group 242: 	165 
    -- CP-element group 242: 	166 
    -- CP-element group 242: 	167 
    -- CP-element group 242: 	168 
    -- CP-element group 242: 	169 
    -- CP-element group 242: 	170 
    -- CP-element group 242: 	176 
    -- CP-element group 242: 	177 
    -- CP-element group 242: 	178 
    -- CP-element group 242: 	179 
    -- CP-element group 242:  members (44) 
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261__entry__
      -- CP-element group 242: 	 branch_block_stmt_785/merge_stmt_1211__exit__
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_update_start_
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_address_calculated
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_root_address_calculated
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_address_resized
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_addr_resize/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_addr_resize/$exit
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_addr_resize/base_resize_req
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_addr_resize/base_resize_ack
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_plus_offset/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_plus_offset/$exit
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_plus_offset/sum_rename_req
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_base_plus_offset/sum_rename_ack
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_sample_start
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_update_start
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_0_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_0_Sample/rr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_0_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_0_Update/cr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_1_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_1_Sample/rr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_1_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_1_Update/cr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_2_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_2_Sample/rr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_2_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_2_Update/cr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_3_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_3_Sample/rr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_3_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_word_addrgen_3_Update/cr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_0/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_0/cr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_1/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_1/cr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_2/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_2/cr
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_3/$entry
      -- CP-element group 242: 	 branch_block_stmt_785/assign_stmt_1247_to_assign_stmt_1261/ptr_deref_1250_Update/word_access_complete/word_3/cr
      -- CP-element group 242: 	 branch_block_stmt_785/merge_stmt_1211_PhiAck/$exit
      -- 
    rr_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_addr_0_req_0); -- 
    cr_4224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_addr_0_req_1); -- 
    rr_4229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_addr_1_req_0); -- 
    cr_4234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_addr_1_req_1); -- 
    rr_4239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_addr_2_req_0); -- 
    cr_4244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_addr_2_req_1); -- 
    rr_4249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_addr_3_req_0); -- 
    cr_4254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_addr_3_req_1); -- 
    cr_4291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_load_0_req_1); -- 
    cr_4296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_load_1_req_1); -- 
    cr_4301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_load_2_req_1); -- 
    cr_4306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(242), ack => ptr_deref_1250_load_3_req_1); -- 
    zeropad3D_A_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_2875_elements(239) & zeropad3D_A_CP_2875_elements(240) & zeropad3D_A_CP_2875_elements(241);
      gj_zeropad3D_A_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_2875_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  merge  transition  place  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	75 
    -- CP-element group 243: 	183 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	184 
    -- CP-element group 243:  members (10) 
      -- CP-element group 243: 	 branch_block_stmt_785/merge_stmt_1270__exit__
      -- CP-element group 243: 	 branch_block_stmt_785/assign_stmt_1274__entry__
      -- CP-element group 243: 	 branch_block_stmt_785/merge_stmt_1270_PhiAck/dummy
      -- CP-element group 243: 	 branch_block_stmt_785/merge_stmt_1270_PhiAck/$exit
      -- CP-element group 243: 	 branch_block_stmt_785/assign_stmt_1274/$entry
      -- CP-element group 243: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_785/merge_stmt_1270_PhiAck/$entry
      -- CP-element group 243: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_785/assign_stmt_1274/WPIPE_Block0_complete_1272_Sample/req
      -- CP-element group 243: 	 branch_block_stmt_785/merge_stmt_1270_PhiReqMerge
      -- 
    req_4342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_2875_elements(243), ack => WPIPE_Block0_complete_1272_inst_req_0); -- 
    zeropad3D_A_CP_2875_elements(243) <= OrReduce(zeropad3D_A_CP_2875_elements(75) & zeropad3D_A_CP_2875_elements(183));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1021_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1100_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1125_wire : std_logic_vector(31 downto 0);
    signal LOAD_pad_791_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_791_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom89_1111_resized : std_logic_vector(13 downto 0);
    signal R_idxprom89_1111_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom94_1136_resized : std_logic_vector(13 downto 0);
    signal R_idxprom94_1136_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1033_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1033_scaled : std_logic_vector(13 downto 0);
    signal add108_1188 : std_logic_vector(31 downto 0);
    signal add122_873 : std_logic_vector(31 downto 0);
    signal add56_1009 : std_logic_vector(31 downto 0);
    signal add60_1014 : std_logic_vector(31 downto 0);
    signal add75_1073 : std_logic_vector(31 downto 0);
    signal add82_1088 : std_logic_vector(31 downto 0);
    signal add86_1093 : std_logic_vector(31 downto 0);
    signal add97_1151 : std_logic_vector(31 downto 0);
    signal add_1256 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1034_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1034_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1034_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1034_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1034_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1034_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1112_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1112_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1112_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1112_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1112_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1112_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1137_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1137_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1137_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1137_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1137_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1137_root_address : std_logic_vector(13 downto 0);
    signal arrayidx90_1114 : std_logic_vector(31 downto 0);
    signal arrayidx95_1139 : std_logic_vector(31 downto 0);
    signal arrayidx_1036 : std_logic_vector(31 downto 0);
    signal call_788 : std_logic_vector(7 downto 0);
    signal cmp100_1158 : std_logic_vector(0 downto 0);
    signal cmp109_1193 : std_logic_vector(0 downto 0);
    signal cmp123_878 : std_logic_vector(0 downto 0);
    signal cmp28_929 : std_logic_vector(0 downto 0);
    signal cmp35x_xnot_946 : std_logic_vector(0 downto 0);
    signal cmp41_953 : std_logic_vector(0 downto 0);
    signal cmp49_987 : std_logic_vector(0 downto 0);
    signal cmp_1261 : std_logic_vector(0 downto 0);
    signal conv_796 : std_logic_vector(31 downto 0);
    signal iNsTr_17_973 : std_logic_vector(31 downto 0);
    signal iNsTr_23_1247 : std_logic_vector(31 downto 0);
    signal iNsTr_25_1179 : std_logic_vector(31 downto 0);
    signal iNsTr_2_804 : std_logic_vector(31 downto 0);
    signal iNsTr_3_816 : std_logic_vector(31 downto 0);
    signal iNsTr_4_828 : std_logic_vector(31 downto 0);
    signal iNsTr_5_840 : std_logic_vector(31 downto 0);
    signal iNsTr_6_857 : std_logic_vector(31 downto 0);
    signal idxprom89_1107 : std_logic_vector(63 downto 0);
    signal idxprom94_1132 : std_logic_vector(63 downto 0);
    signal idxprom_1029 : std_logic_vector(63 downto 0);
    signal inc114_1197 : std_logic_vector(31 downto 0);
    signal inc114x_xix_x1_1202 : std_logic_vector(31 downto 0);
    signal inc_1171 : std_logic_vector(31 downto 0);
    signal ix_x0_1231 : std_logic_vector(31 downto 0);
    signal ix_x1126_900 : std_logic_vector(31 downto 0);
    signal jx_x0_1212 : std_logic_vector(31 downto 0);
    signal jx_x1124_914 : std_logic_vector(31 downto 0);
    signal kx_x0125_907 : std_logic_vector(31 downto 0);
    signal kx_x1_1221 : std_logic_vector(31 downto 0);
    signal mul19_849 : std_logic_vector(31 downto 0);
    signal mul24121_867 : std_logic_vector(31 downto 0);
    signal mul55_999 : std_logic_vector(31 downto 0);
    signal mul59_1004 : std_logic_vector(31 downto 0);
    signal mul74_1058 : std_logic_vector(31 downto 0);
    signal mul81_1078 : std_logic_vector(31 downto 0);
    signal mul85_1083 : std_logic_vector(31 downto 0);
    signal orx_xcond_958 : std_logic_vector(0 downto 0);
    signal ptr_deref_1038_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1038_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1038_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1038_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1038_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1038_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1117_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1117_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1117_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1117_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1117_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1141_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1141_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1141_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1141_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1141_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1141_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1182_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1182_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1182_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1182_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1182_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_1182_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1250_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1250_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1250_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1250_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_1250_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_807_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_807_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_807_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_807_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_807_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_807_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_807_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_807_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_807_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_807_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_807_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_807_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_807_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_807_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_819_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_819_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_819_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_819_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_819_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_819_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_819_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_819_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_819_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_819_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_819_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_819_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_819_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_819_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_831_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_831_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_831_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_831_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_831_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_843_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_843_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_843_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_843_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_843_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_860_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_860_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_860_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_860_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_860_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_860_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_860_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_860_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_860_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_860_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_860_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_860_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_860_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_860_word_offset_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_976_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_976_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_976_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_976_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_976_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_976_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_976_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_976_word_address_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_976_word_address_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_976_word_address_3 : std_logic_vector(8 downto 0);
    signal ptr_deref_976_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_976_word_offset_1 : std_logic_vector(8 downto 0);
    signal ptr_deref_976_word_offset_2 : std_logic_vector(8 downto 0);
    signal ptr_deref_976_word_offset_3 : std_logic_vector(8 downto 0);
    signal shr88_1102 : std_logic_vector(31 downto 0);
    signal shr93_1127 : std_logic_vector(31 downto 0);
    signal shr_1023 : std_logic_vector(31 downto 0);
    signal sub34_941 : std_logic_vector(31 downto 0);
    signal sub48_982 : std_logic_vector(31 downto 0);
    signal sub67_1048 : std_logic_vector(31 downto 0);
    signal sub73_1053 : std_logic_vector(31 downto 0);
    signal sub_891 : std_logic_vector(31 downto 0);
    signal tmp105_1183 : std_logic_vector(31 downto 0);
    signal tmp10_844 : std_logic_vector(31 downto 0);
    signal tmp118_1063 : std_logic_vector(31 downto 0);
    signal tmp119_1068 : std_logic_vector(31 downto 0);
    signal tmp22120_861 : std_logic_vector(31 downto 0);
    signal tmp22_1251 : std_logic_vector(31 downto 0);
    signal tmp2_808 : std_logic_vector(31 downto 0);
    signal tmp31_894 : std_logic_vector(31 downto 0);
    signal tmp45_977 : std_logic_vector(31 downto 0);
    signal tmp4_820 : std_logic_vector(31 downto 0);
    signal tmp8_832 : std_logic_vector(31 downto 0);
    signal tmp91_1118 : std_logic_vector(63 downto 0);
    signal tmp_792 : std_logic_vector(7 downto 0);
    signal type_cast_1017_wire : std_logic_vector(31 downto 0);
    signal type_cast_1020_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1027_wire : std_logic_vector(63 downto 0);
    signal type_cast_1040_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1096_wire : std_logic_vector(31 downto 0);
    signal type_cast_1099_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1105_wire : std_logic_vector(63 downto 0);
    signal type_cast_1121_wire : std_logic_vector(31 downto 0);
    signal type_cast_1124_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1130_wire : std_logic_vector(63 downto 0);
    signal type_cast_1149_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1154_wire : std_logic_vector(31 downto 0);
    signal type_cast_1156_wire : std_logic_vector(31 downto 0);
    signal type_cast_1169_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1216_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1218_wire : std_logic_vector(31 downto 0);
    signal type_cast_1220_wire : std_logic_vector(31 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1228_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1230_wire : std_logic_vector(31 downto 0);
    signal type_cast_1234_wire : std_logic_vector(31 downto 0);
    signal type_cast_1236_wire : std_logic_vector(31 downto 0);
    signal type_cast_1238_wire : std_logic_vector(31 downto 0);
    signal type_cast_865_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_870_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_889_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_897_wire : std_logic_vector(31 downto 0);
    signal type_cast_899_wire : std_logic_vector(31 downto 0);
    signal type_cast_904_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_906_wire : std_logic_vector(31 downto 0);
    signal type_cast_911_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_913_wire : std_logic_vector(31 downto 0);
    signal type_cast_918_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_920_wire : std_logic_vector(31 downto 0);
    signal type_cast_925_wire : std_logic_vector(31 downto 0);
    signal type_cast_927_wire : std_logic_vector(31 downto 0);
    signal type_cast_949_wire : std_logic_vector(31 downto 0);
    signal type_cast_951_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_pad_791_word_address_0 <= "0";
    array_obj_ref_1034_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1034_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1034_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1034_resized_base_address <= "00000000000000";
    array_obj_ref_1112_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1112_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1112_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1112_resized_base_address <= "00000000000000";
    array_obj_ref_1137_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1137_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1137_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1137_resized_base_address <= "00000000000000";
    iNsTr_17_973 <= "00000000000000000000000000001101";
    iNsTr_23_1247 <= "00000000000000000000000000001001";
    iNsTr_25_1179 <= "00000000000000000000000000001101";
    iNsTr_2_804 <= "00000000000000000000000000010001";
    iNsTr_3_816 <= "00000000000000000000000000001101";
    iNsTr_4_828 <= "00000000000000000000000000000100";
    iNsTr_5_840 <= "00000000000000000000000000000011";
    iNsTr_6_857 <= "00000000000000000000000000001001";
    ptr_deref_1038_word_offset_0 <= "00000000000000";
    ptr_deref_1117_word_offset_0 <= "00000000000000";
    ptr_deref_1141_word_offset_0 <= "00000000000000";
    ptr_deref_1182_word_offset_0 <= "000000000";
    ptr_deref_1182_word_offset_1 <= "000000001";
    ptr_deref_1182_word_offset_2 <= "000000010";
    ptr_deref_1182_word_offset_3 <= "000000011";
    ptr_deref_1250_word_offset_0 <= "000000000";
    ptr_deref_1250_word_offset_1 <= "000000001";
    ptr_deref_1250_word_offset_2 <= "000000010";
    ptr_deref_1250_word_offset_3 <= "000000011";
    ptr_deref_807_word_offset_0 <= "000000000";
    ptr_deref_807_word_offset_1 <= "000000001";
    ptr_deref_807_word_offset_2 <= "000000010";
    ptr_deref_807_word_offset_3 <= "000000011";
    ptr_deref_819_word_offset_0 <= "000000000";
    ptr_deref_819_word_offset_1 <= "000000001";
    ptr_deref_819_word_offset_2 <= "000000010";
    ptr_deref_819_word_offset_3 <= "000000011";
    ptr_deref_831_word_offset_0 <= "0000000";
    ptr_deref_843_word_offset_0 <= "0000000";
    ptr_deref_860_word_offset_0 <= "000000000";
    ptr_deref_860_word_offset_1 <= "000000001";
    ptr_deref_860_word_offset_2 <= "000000010";
    ptr_deref_860_word_offset_3 <= "000000011";
    ptr_deref_976_word_offset_0 <= "000000000";
    ptr_deref_976_word_offset_1 <= "000000001";
    ptr_deref_976_word_offset_2 <= "000000010";
    ptr_deref_976_word_offset_3 <= "000000011";
    type_cast_1020_wire_constant <= "00000000000000000000000000000010";
    type_cast_1040_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1099_wire_constant <= "00000000000000000000000000000010";
    type_cast_1124_wire_constant <= "00000000000000000000000000000010";
    type_cast_1149_wire_constant <= "00000000000000000000000000000100";
    type_cast_1169_wire_constant <= "00000000000000000000000000000001";
    type_cast_1216_wire_constant <= "00000000000000000000000000000000";
    type_cast_1225_wire_constant <= "00000000000000000000000000000000";
    type_cast_1228_wire_constant <= "00000000000000000000000000000000";
    type_cast_865_wire_constant <= "00000000000000000000000000000001";
    type_cast_870_wire_constant <= "00000000000000000000000000000000";
    type_cast_889_wire_constant <= "11111111111111111111111111111111";
    type_cast_904_wire_constant <= "00000000000000000000000000000000";
    type_cast_911_wire_constant <= "00000000000000000000000000000000";
    type_cast_918_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_1212: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_1216_wire_constant & type_cast_1218_wire & type_cast_1220_wire;
      req <= phi_stmt_1212_req_0 & phi_stmt_1212_req_1 & phi_stmt_1212_req_2;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1212",
          num_reqs => 3,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1212_ack_0,
          idata => idata,
          odata => jx_x0_1212,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1212
    phi_stmt_1221: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_1225_wire_constant & type_cast_1228_wire_constant & type_cast_1230_wire;
      req <= phi_stmt_1221_req_0 & phi_stmt_1221_req_1 & phi_stmt_1221_req_2;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1221",
          num_reqs => 3,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1221_ack_0,
          idata => idata,
          odata => kx_x1_1221,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1221
    phi_stmt_1231: Block -- phi operator 
      signal idata: std_logic_vector(95 downto 0);
      signal req: BooleanArray(2 downto 0);
      --
    begin -- 
      idata <= type_cast_1234_wire & type_cast_1236_wire & type_cast_1238_wire;
      req <= phi_stmt_1231_req_0 & phi_stmt_1231_req_1 & phi_stmt_1231_req_2;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1231",
          num_reqs => 3,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1231_ack_0,
          idata => idata,
          odata => ix_x0_1231,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1231
    phi_stmt_894: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_897_wire & type_cast_899_wire;
      req <= phi_stmt_894_req_0 & phi_stmt_894_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_894",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_894_ack_0,
          idata => idata,
          odata => tmp31_894,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_894
    phi_stmt_900: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_904_wire_constant & type_cast_906_wire;
      req <= phi_stmt_900_req_0 & phi_stmt_900_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_900",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_900_ack_0,
          idata => idata,
          odata => ix_x1126_900,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_900
    phi_stmt_907: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_911_wire_constant & type_cast_913_wire;
      req <= phi_stmt_907_req_0 & phi_stmt_907_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_907",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_907_ack_0,
          idata => idata,
          odata => kx_x0125_907,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_907
    phi_stmt_914: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_918_wire_constant & type_cast_920_wire;
      req <= phi_stmt_914_req_0 & phi_stmt_914_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_914",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_914_ack_0,
          idata => idata,
          odata => jx_x1124_914,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_914
    addr_of_1035_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1035_final_reg_req_0;
      addr_of_1035_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1035_final_reg_req_1;
      addr_of_1035_final_reg_ack_1<= rack(0);
      addr_of_1035_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1035_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1034_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1036,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1113_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1113_final_reg_req_0;
      addr_of_1113_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1113_final_reg_req_1;
      addr_of_1113_final_reg_ack_1<= rack(0);
      addr_of_1113_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1113_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1112_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx90_1114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1138_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1138_final_reg_req_0;
      addr_of_1138_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1138_final_reg_req_1;
      addr_of_1138_final_reg_ack_1<= rack(0);
      addr_of_1138_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1138_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1137_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx95_1139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1017_inst
    process(add60_1014) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add60_1014(31 downto 0);
      type_cast_1017_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1022_inst
    process(ASHR_i32_i32_1021_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1021_wire(31 downto 0);
      shr_1023 <= tmp_var; -- 
    end process;
    type_cast_1028_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1028_inst_req_0;
      type_cast_1028_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1028_inst_req_1;
      type_cast_1028_inst_ack_1<= rack(0);
      type_cast_1028_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1028_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1027_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1029,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1096_inst
    process(add75_1073) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add75_1073(31 downto 0);
      type_cast_1096_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1101_inst
    process(ASHR_i32_i32_1100_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1100_wire(31 downto 0);
      shr88_1102 <= tmp_var; -- 
    end process;
    type_cast_1106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1106_inst_req_0;
      type_cast_1106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1106_inst_req_1;
      type_cast_1106_inst_ack_1<= rack(0);
      type_cast_1106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1105_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom89_1107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1121_inst
    process(add86_1093) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add86_1093(31 downto 0);
      type_cast_1121_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1126_inst
    process(ASHR_i32_i32_1125_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1125_wire(31 downto 0);
      shr93_1127 <= tmp_var; -- 
    end process;
    type_cast_1131_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1131_inst_req_0;
      type_cast_1131_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1131_inst_req_1;
      type_cast_1131_inst_ack_1<= rack(0);
      type_cast_1131_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1131_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1130_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom94_1132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1154_inst
    process(add97_1151) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add97_1151(31 downto 0);
      type_cast_1154_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1156_inst
    process(tmp2_808) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := tmp2_808(31 downto 0);
      type_cast_1156_wire <= tmp_var; -- 
    end process;
    type_cast_1196_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1196_inst_req_0;
      type_cast_1196_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1196_inst_req_1;
      type_cast_1196_inst_ack_1<= rack(0);
      type_cast_1196_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1196_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp109_1193,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc114_1197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1218_inst_req_0;
      type_cast_1218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1218_inst_req_1;
      type_cast_1218_inst_ack_1<= rack(0);
      type_cast_1218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1218_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1220_inst_req_0;
      type_cast_1220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1220_inst_req_1;
      type_cast_1220_inst_ack_1<= rack(0);
      type_cast_1220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1124_914,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1220_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1230_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1230_inst_req_0;
      type_cast_1230_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1230_inst_req_1;
      type_cast_1230_inst_ack_1<= rack(0);
      type_cast_1230_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1230_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add97_1151,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1230_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1234_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1234_inst_req_0;
      type_cast_1234_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1234_inst_req_1;
      type_cast_1234_inst_ack_1<= rack(0);
      type_cast_1234_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1234_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc114x_xix_x1_1202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1234_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1236_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1236_inst_req_0;
      type_cast_1236_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1236_inst_req_1;
      type_cast_1236_inst_ack_1<= rack(0);
      type_cast_1236_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1236_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc114x_xix_x1_1202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1236_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1126_900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1238_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_795_inst_req_0;
      type_cast_795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_795_inst_req_1;
      type_cast_795_inst_ack_1<= rack(0);
      type_cast_795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_897_inst_req_0;
      type_cast_897_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_897_inst_req_1;
      type_cast_897_inst_ack_1<= rack(0);
      type_cast_897_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_897_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp22120_861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_897_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_899_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_899_inst_req_0;
      type_cast_899_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_899_inst_req_1;
      type_cast_899_inst_ack_1<= rack(0);
      type_cast_899_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_899_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp22_1251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_899_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_906_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_906_inst_req_0;
      type_cast_906_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_906_inst_req_1;
      type_cast_906_inst_ack_1<= rack(0);
      type_cast_906_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_906_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x0_1231,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_906_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_913_inst_req_0;
      type_cast_913_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_913_inst_req_1;
      type_cast_913_inst_ack_1<= rack(0);
      type_cast_913_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_913_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x1_1221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_913_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_920_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_920_inst_req_0;
      type_cast_920_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_920_inst_req_1;
      type_cast_920_inst_ack_1<= rack(0);
      type_cast_920_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_920_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0_1212,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_920_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_925_inst
    process(ix_x1126_900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ix_x1126_900(31 downto 0);
      type_cast_925_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_927_inst
    process(sub_891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sub_891(31 downto 0);
      type_cast_927_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_949_inst
    process(jx_x1124_914) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := jx_x1124_914(31 downto 0);
      type_cast_949_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_951_inst
    process(sub_891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sub_891(31 downto 0);
      type_cast_951_wire <= tmp_var; -- 
    end process;
    -- equivalence LOAD_pad_791_gather_scatter
    process(LOAD_pad_791_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_791_data_0;
      ov(7 downto 0) := iv;
      tmp_792 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1034_index_1_rename
    process(R_idxprom_1033_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1033_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1033_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1034_index_1_resize
    process(idxprom_1029) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1029;
      ov := iv(13 downto 0);
      R_idxprom_1033_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1034_root_address_inst
    process(array_obj_ref_1034_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1034_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1034_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1112_index_1_rename
    process(R_idxprom89_1111_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom89_1111_resized;
      ov(13 downto 0) := iv;
      R_idxprom89_1111_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1112_index_1_resize
    process(idxprom89_1107) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom89_1107;
      ov := iv(13 downto 0);
      R_idxprom89_1111_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1112_root_address_inst
    process(array_obj_ref_1112_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1112_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1112_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1137_index_1_rename
    process(R_idxprom94_1136_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom94_1136_resized;
      ov(13 downto 0) := iv;
      R_idxprom94_1136_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1137_index_1_resize
    process(idxprom94_1132) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom94_1132;
      ov := iv(13 downto 0);
      R_idxprom94_1136_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1137_root_address_inst
    process(array_obj_ref_1137_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1137_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1137_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1038_addr_0
    process(ptr_deref_1038_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1038_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1038_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1038_base_resize
    process(arrayidx_1036) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1036;
      ov := iv(13 downto 0);
      ptr_deref_1038_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1038_gather_scatter
    process(type_cast_1040_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1040_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1038_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1038_root_address_inst
    process(ptr_deref_1038_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1038_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1038_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1117_addr_0
    process(ptr_deref_1117_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1117_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1117_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1117_base_resize
    process(arrayidx90_1114) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx90_1114;
      ov := iv(13 downto 0);
      ptr_deref_1117_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1117_gather_scatter
    process(ptr_deref_1117_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1117_data_0;
      ov(63 downto 0) := iv;
      tmp91_1118 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1117_root_address_inst
    process(ptr_deref_1117_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1117_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1117_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1141_addr_0
    process(ptr_deref_1141_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1141_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1141_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1141_base_resize
    process(arrayidx95_1139) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx95_1139;
      ov := iv(13 downto 0);
      ptr_deref_1141_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1141_gather_scatter
    process(tmp91_1118) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp91_1118;
      ov(63 downto 0) := iv;
      ptr_deref_1141_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1141_root_address_inst
    process(ptr_deref_1141_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1141_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1141_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1182_base_resize
    process(iNsTr_25_1179) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_25_1179;
      ov := iv(8 downto 0);
      ptr_deref_1182_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1182_gather_scatter
    process(ptr_deref_1182_data_3, ptr_deref_1182_data_2, ptr_deref_1182_data_1, ptr_deref_1182_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1182_data_3 & ptr_deref_1182_data_2 & ptr_deref_1182_data_1 & ptr_deref_1182_data_0;
      ov(31 downto 0) := iv;
      tmp105_1183 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1182_root_address_inst
    process(ptr_deref_1182_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1182_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_1182_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1250_base_resize
    process(iNsTr_23_1247) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_23_1247;
      ov := iv(8 downto 0);
      ptr_deref_1250_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1250_gather_scatter
    process(ptr_deref_1250_data_3, ptr_deref_1250_data_2, ptr_deref_1250_data_1, ptr_deref_1250_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1250_data_3 & ptr_deref_1250_data_2 & ptr_deref_1250_data_1 & ptr_deref_1250_data_0;
      ov(31 downto 0) := iv;
      tmp22_1251 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1250_root_address_inst
    process(ptr_deref_1250_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1250_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_1250_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_807_base_resize
    process(iNsTr_2_804) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_804;
      ov := iv(8 downto 0);
      ptr_deref_807_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_807_gather_scatter
    process(ptr_deref_807_data_3, ptr_deref_807_data_2, ptr_deref_807_data_1, ptr_deref_807_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_807_data_3 & ptr_deref_807_data_2 & ptr_deref_807_data_1 & ptr_deref_807_data_0;
      ov(31 downto 0) := iv;
      tmp2_808 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_807_root_address_inst
    process(ptr_deref_807_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_807_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_807_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_819_base_resize
    process(iNsTr_3_816) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_816;
      ov := iv(8 downto 0);
      ptr_deref_819_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_819_gather_scatter
    process(ptr_deref_819_data_3, ptr_deref_819_data_2, ptr_deref_819_data_1, ptr_deref_819_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_819_data_3 & ptr_deref_819_data_2 & ptr_deref_819_data_1 & ptr_deref_819_data_0;
      ov(31 downto 0) := iv;
      tmp4_820 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_819_root_address_inst
    process(ptr_deref_819_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_819_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_819_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_831_addr_0
    process(ptr_deref_831_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_831_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_831_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_831_base_resize
    process(iNsTr_4_828) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_828;
      ov := iv(6 downto 0);
      ptr_deref_831_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_831_gather_scatter
    process(ptr_deref_831_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_831_data_0;
      ov(31 downto 0) := iv;
      tmp8_832 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_831_root_address_inst
    process(ptr_deref_831_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_831_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_831_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_843_addr_0
    process(ptr_deref_843_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_843_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_843_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_843_base_resize
    process(iNsTr_5_840) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_840;
      ov := iv(6 downto 0);
      ptr_deref_843_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_843_gather_scatter
    process(ptr_deref_843_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_843_data_0;
      ov(31 downto 0) := iv;
      tmp10_844 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_843_root_address_inst
    process(ptr_deref_843_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_843_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_843_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_860_base_resize
    process(iNsTr_6_857) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_857;
      ov := iv(8 downto 0);
      ptr_deref_860_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_860_gather_scatter
    process(ptr_deref_860_data_3, ptr_deref_860_data_2, ptr_deref_860_data_1, ptr_deref_860_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_860_data_3 & ptr_deref_860_data_2 & ptr_deref_860_data_1 & ptr_deref_860_data_0;
      ov(31 downto 0) := iv;
      tmp22120_861 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_860_root_address_inst
    process(ptr_deref_860_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_860_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_860_root_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_976_base_resize
    process(iNsTr_17_973) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_973;
      ov := iv(8 downto 0);
      ptr_deref_976_resized_base_address <= ov(8 downto 0);
      --
    end process;
    -- equivalence ptr_deref_976_gather_scatter
    process(ptr_deref_976_data_3, ptr_deref_976_data_2, ptr_deref_976_data_1, ptr_deref_976_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_976_data_3 & ptr_deref_976_data_2 & ptr_deref_976_data_1 & ptr_deref_976_data_0;
      ov(31 downto 0) := iv;
      tmp45_977 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_976_root_address_inst
    process(ptr_deref_976_resized_base_address) --
      variable iv : std_logic_vector(8 downto 0);
      variable ov : std_logic_vector(8 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_976_resized_base_address;
      ov(8 downto 0) := iv;
      ptr_deref_976_root_address <= ov(8 downto 0);
      --
    end process;
    if_stmt_1159_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp100_1158;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1159_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1159_branch_req_0,
          ack0 => if_stmt_1159_branch_ack_0,
          ack1 => if_stmt_1159_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1203_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp109_1193;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1203_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1203_branch_req_0,
          ack0 => if_stmt_1203_branch_ack_0,
          ack1 => if_stmt_1203_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1262_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1261;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1262_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1262_branch_req_0,
          ack0 => if_stmt_1262_branch_ack_0,
          ack1 => if_stmt_1262_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_879_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp123_878;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_879_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_879_branch_req_0,
          ack0 => if_stmt_879_branch_ack_0,
          ack1 => if_stmt_879_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_930_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp28_929;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_930_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_930_branch_req_0,
          ack0 => if_stmt_930_branch_ack_0,
          ack1 => if_stmt_930_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_959_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_958;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_959_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_959_branch_req_0,
          ack0 => if_stmt_959_branch_ack_0,
          ack1 => if_stmt_959_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_988_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp49_987;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_988_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_988_branch_req_0,
          ack0 => if_stmt_988_branch_ack_0,
          ack1 => if_stmt_988_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1008_inst
    process(kx_x0125_907, mul55_999) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x0125_907, mul55_999, tmp_var);
      add56_1009 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1013_inst
    process(add56_1009, mul59_1004) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add56_1009, mul59_1004, tmp_var);
      add60_1014 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1062_inst
    process(mul74_1058, sub67_1048) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1058, sub67_1048, tmp_var);
      tmp118_1063 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1072_inst
    process(tmp119_1068, kx_x0125_907) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp119_1068, kx_x0125_907, tmp_var);
      add75_1073 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1087_inst
    process(kx_x0125_907, mul81_1078) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x0125_907, mul81_1078, tmp_var);
      add82_1088 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1092_inst
    process(add82_1088, mul85_1083) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add82_1088, mul85_1083, tmp_var);
      add86_1093 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1150_inst
    process(kx_x0125_907) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x0125_907, type_cast_1149_wire_constant, tmp_var);
      add97_1151 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1170_inst
    process(jx_x1124_914) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1124_914, type_cast_1169_wire_constant, tmp_var);
      inc_1171 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1187_inst
    process(tmp105_1183, mul24121_867) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp105_1183, mul24121_867, tmp_var);
      add108_1188 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1201_inst
    process(inc114_1197, ix_x1126_900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc114_1197, ix_x1126_900, tmp_var);
      inc114x_xix_x1_1202 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1255_inst
    process(tmp22_1251, mul24121_867) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp22_1251, mul24121_867, tmp_var);
      add_1256 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_890_inst
    process(conv_796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv_796, type_cast_889_wire_constant, tmp_var);
      sub_891 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_940_inst
    process(sub_891, tmp31_894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_891, tmp31_894, tmp_var);
      sub34_941 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_981_inst
    process(sub_891, tmp45_977) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_891, tmp45_977, tmp_var);
      sub48_982 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_957_inst
    process(cmp35x_xnot_946, cmp41_953) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp35x_xnot_946, cmp41_953, tmp_var);
      orx_xcond_958 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1021_inst
    process(type_cast_1017_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1017_wire, type_cast_1020_wire_constant, tmp_var);
      ASHR_i32_i32_1021_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1100_inst
    process(type_cast_1096_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1096_wire, type_cast_1099_wire_constant, tmp_var);
      ASHR_i32_i32_1100_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1125_inst
    process(type_cast_1121_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1121_wire, type_cast_1124_wire_constant, tmp_var);
      ASHR_i32_i32_1125_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1192_inst
    process(inc_1171, add108_1188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1171, add108_1188, tmp_var);
      cmp109_1193 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_877_inst
    process(tmp22120_861, add122_873) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tmp22120_861, add122_873, tmp_var);
      cmp123_878 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1003_inst
    process(ix_x1126_900, mul19_849) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(ix_x1126_900, mul19_849, tmp_var);
      mul59_1004 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1057_inst
    process(tmp4_820, sub73_1053) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp4_820, sub73_1053, tmp_var);
      mul74_1058 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1067_inst
    process(tmp118_1063, tmp2_808) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp118_1063, tmp2_808, tmp_var);
      tmp119_1068 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1077_inst
    process(jx_x1124_914, tmp8_832) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(jx_x1124_914, tmp8_832, tmp_var);
      mul81_1078 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1082_inst
    process(ix_x1126_900, mul19_849) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(ix_x1126_900, mul19_849, tmp_var);
      mul85_1083 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_848_inst
    process(tmp10_844, tmp8_832) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp10_844, tmp8_832, tmp_var);
      mul19_849 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_998_inst
    process(jx_x1124_914, tmp8_832) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(jx_x1124_914, tmp8_832, tmp_var);
      mul55_999 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_928_inst
    process(type_cast_925_wire, type_cast_927_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_925_wire, type_cast_927_wire, tmp_var);
      cmp28_929 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_952_inst
    process(type_cast_949_wire, type_cast_951_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_949_wire, type_cast_951_wire, tmp_var);
      cmp41_953 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_866_inst
    process(conv_796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_796, type_cast_865_wire_constant, tmp_var);
      mul24121_867 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1157_inst
    process(type_cast_1154_wire, type_cast_1156_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1154_wire, type_cast_1156_wire, tmp_var);
      cmp100_1158 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1047_inst
    process(jx_x1124_914, conv_796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(jx_x1124_914, conv_796, tmp_var);
      sub67_1048 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1052_inst
    process(ix_x1126_900, conv_796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(ix_x1126_900, conv_796, tmp_var);
      sub73_1053 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_872_inst
    process(type_cast_870_wire_constant, mul24121_867) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(type_cast_870_wire_constant, mul24121_867, tmp_var);
      add122_873 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_986_inst
    process(jx_x1124_914, sub48_982) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(jx_x1124_914, sub48_982, tmp_var);
      cmp49_987 <= tmp_var; --
    end process;
    -- binary operator ULE_u32_u1_945_inst
    process(ix_x1126_900, sub34_941) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(ix_x1126_900, sub34_941, tmp_var);
      cmp35x_xnot_946 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1260_inst
    process(ix_x0_1231, add_1256) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(ix_x0_1231, add_1256, tmp_var);
      cmp_1261 <= tmp_var; --
    end process;
    -- shared split operator group (37) : array_obj_ref_1034_index_offset 
    ApIntAdd_group_37: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1033_scaled;
      array_obj_ref_1034_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1034_index_offset_req_0;
      array_obj_ref_1034_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1034_index_offset_req_1;
      array_obj_ref_1034_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_37_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : array_obj_ref_1112_index_offset 
    ApIntAdd_group_38: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom89_1111_scaled;
      array_obj_ref_1112_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1112_index_offset_req_0;
      array_obj_ref_1112_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1112_index_offset_req_1;
      array_obj_ref_1112_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_38_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : array_obj_ref_1137_index_offset 
    ApIntAdd_group_39: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom94_1136_scaled;
      array_obj_ref_1137_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1137_index_offset_req_0;
      array_obj_ref_1137_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1137_index_offset_req_1;
      array_obj_ref_1137_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_39_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_39_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : ptr_deref_1182_addr_0 
    ApIntAdd_group_40: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1182_root_address;
      ptr_deref_1182_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1182_addr_0_req_0;
      ptr_deref_1182_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1182_addr_0_req_1;
      ptr_deref_1182_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_40_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_40_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_40",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : ptr_deref_1182_addr_1 
    ApIntAdd_group_41: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1182_root_address;
      ptr_deref_1182_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1182_addr_1_req_0;
      ptr_deref_1182_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1182_addr_1_req_1;
      ptr_deref_1182_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_41_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_41_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : ptr_deref_1182_addr_2 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1182_root_address;
      ptr_deref_1182_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1182_addr_2_req_0;
      ptr_deref_1182_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1182_addr_2_req_1;
      ptr_deref_1182_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : ptr_deref_1182_addr_3 
    ApIntAdd_group_43: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1182_root_address;
      ptr_deref_1182_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1182_addr_3_req_0;
      ptr_deref_1182_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1182_addr_3_req_1;
      ptr_deref_1182_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_43_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_43_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_43",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : ptr_deref_1250_addr_0 
    ApIntAdd_group_44: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1250_root_address;
      ptr_deref_1250_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1250_addr_0_req_0;
      ptr_deref_1250_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1250_addr_0_req_1;
      ptr_deref_1250_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_44_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_44_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : ptr_deref_1250_addr_1 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1250_root_address;
      ptr_deref_1250_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1250_addr_1_req_0;
      ptr_deref_1250_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1250_addr_1_req_1;
      ptr_deref_1250_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : ptr_deref_1250_addr_2 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1250_root_address;
      ptr_deref_1250_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1250_addr_2_req_0;
      ptr_deref_1250_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1250_addr_2_req_1;
      ptr_deref_1250_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : ptr_deref_1250_addr_3 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_1250_root_address;
      ptr_deref_1250_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_1250_addr_3_req_0;
      ptr_deref_1250_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1250_addr_3_req_1;
      ptr_deref_1250_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : ptr_deref_807_addr_0 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_807_root_address;
      ptr_deref_807_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_807_addr_0_req_0;
      ptr_deref_807_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_807_addr_0_req_1;
      ptr_deref_807_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : ptr_deref_807_addr_1 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_807_root_address;
      ptr_deref_807_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_807_addr_1_req_0;
      ptr_deref_807_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_807_addr_1_req_1;
      ptr_deref_807_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : ptr_deref_807_addr_2 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_807_root_address;
      ptr_deref_807_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_807_addr_2_req_0;
      ptr_deref_807_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_807_addr_2_req_1;
      ptr_deref_807_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : ptr_deref_807_addr_3 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_807_root_address;
      ptr_deref_807_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_807_addr_3_req_0;
      ptr_deref_807_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_807_addr_3_req_1;
      ptr_deref_807_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : ptr_deref_819_addr_0 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_819_root_address;
      ptr_deref_819_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_819_addr_0_req_0;
      ptr_deref_819_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_819_addr_0_req_1;
      ptr_deref_819_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : ptr_deref_819_addr_1 
    ApIntAdd_group_53: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_819_root_address;
      ptr_deref_819_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_819_addr_1_req_0;
      ptr_deref_819_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_819_addr_1_req_1;
      ptr_deref_819_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_53_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_53_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : ptr_deref_819_addr_2 
    ApIntAdd_group_54: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_819_root_address;
      ptr_deref_819_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_819_addr_2_req_0;
      ptr_deref_819_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_819_addr_2_req_1;
      ptr_deref_819_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_54_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_54_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_54",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : ptr_deref_819_addr_3 
    ApIntAdd_group_55: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_819_root_address;
      ptr_deref_819_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_819_addr_3_req_0;
      ptr_deref_819_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_819_addr_3_req_1;
      ptr_deref_819_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_55_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_55_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_55",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : ptr_deref_860_addr_0 
    ApIntAdd_group_56: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_860_root_address;
      ptr_deref_860_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_860_addr_0_req_0;
      ptr_deref_860_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_860_addr_0_req_1;
      ptr_deref_860_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_56_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_56_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_56",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : ptr_deref_860_addr_1 
    ApIntAdd_group_57: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_860_root_address;
      ptr_deref_860_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_860_addr_1_req_0;
      ptr_deref_860_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_860_addr_1_req_1;
      ptr_deref_860_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_57_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_57_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_57",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : ptr_deref_860_addr_2 
    ApIntAdd_group_58: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_860_root_address;
      ptr_deref_860_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_860_addr_2_req_0;
      ptr_deref_860_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_860_addr_2_req_1;
      ptr_deref_860_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_58_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_58_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_58",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : ptr_deref_860_addr_3 
    ApIntAdd_group_59: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_860_root_address;
      ptr_deref_860_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_860_addr_3_req_0;
      ptr_deref_860_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_860_addr_3_req_1;
      ptr_deref_860_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_59_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_59_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_59",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : ptr_deref_976_addr_0 
    ApIntAdd_group_60: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_976_root_address;
      ptr_deref_976_word_address_0 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_976_addr_0_req_0;
      ptr_deref_976_addr_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_976_addr_0_req_1;
      ptr_deref_976_addr_0_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_60_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_60_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : ptr_deref_976_addr_1 
    ApIntAdd_group_61: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_976_root_address;
      ptr_deref_976_word_address_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_976_addr_1_req_0;
      ptr_deref_976_addr_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_976_addr_1_req_1;
      ptr_deref_976_addr_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_61_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_61_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_61",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000001",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : ptr_deref_976_addr_2 
    ApIntAdd_group_62: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_976_root_address;
      ptr_deref_976_word_address_2 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_976_addr_2_req_0;
      ptr_deref_976_addr_2_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_976_addr_2_req_1;
      ptr_deref_976_addr_2_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_62_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_62_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_62",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000010",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : ptr_deref_976_addr_3 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ptr_deref_976_root_address;
      ptr_deref_976_word_address_3 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ptr_deref_976_addr_3_req_0;
      ptr_deref_976_addr_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_976_addr_3_req_1;
      ptr_deref_976_addr_3_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_63_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_63_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000011",
          constant_width => 9,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- unary operator type_cast_1027_inst
    process(shr_1023) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1023, tmp_var);
      type_cast_1027_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1105_inst
    process(shr88_1102) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr88_1102, tmp_var);
      type_cast_1105_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1130_inst
    process(shr93_1127) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr93_1127, tmp_var);
      type_cast_1130_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_pad_791_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_pad_791_load_0_req_0;
      LOAD_pad_791_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_pad_791_load_0_req_1;
      LOAD_pad_791_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_791_word_address_0;
      LOAD_pad_791_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(7 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1117_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1117_load_0_req_0;
      ptr_deref_1117_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1117_load_0_req_1;
      ptr_deref_1117_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1117_word_address_0;
      ptr_deref_1117_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_819_load_3 ptr_deref_807_load_1 ptr_deref_819_load_2 ptr_deref_860_load_3 ptr_deref_860_load_1 ptr_deref_819_load_0 ptr_deref_807_load_0 ptr_deref_860_load_0 ptr_deref_860_load_2 ptr_deref_819_load_1 ptr_deref_807_load_2 ptr_deref_807_load_3 ptr_deref_976_load_0 ptr_deref_976_load_1 ptr_deref_976_load_2 ptr_deref_976_load_3 ptr_deref_1182_load_0 ptr_deref_1182_load_1 ptr_deref_1182_load_2 ptr_deref_1182_load_3 ptr_deref_1250_load_0 ptr_deref_1250_load_1 ptr_deref_1250_load_2 ptr_deref_1250_load_3 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(215 downto 0);
      signal data_out: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 23 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 23 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 23 downto 0);
      signal guard_vector : std_logic_vector( 23 downto 0);
      constant inBUFs : IntegerArray(23 downto 0) := (23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(23 downto 0) := (23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(23 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false);
      constant guardBuffering: IntegerArray(23 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2);
      -- 
    begin -- 
      reqL_unguarded(23) <= ptr_deref_819_load_3_req_0;
      reqL_unguarded(22) <= ptr_deref_807_load_1_req_0;
      reqL_unguarded(21) <= ptr_deref_819_load_2_req_0;
      reqL_unguarded(20) <= ptr_deref_860_load_3_req_0;
      reqL_unguarded(19) <= ptr_deref_860_load_1_req_0;
      reqL_unguarded(18) <= ptr_deref_819_load_0_req_0;
      reqL_unguarded(17) <= ptr_deref_807_load_0_req_0;
      reqL_unguarded(16) <= ptr_deref_860_load_0_req_0;
      reqL_unguarded(15) <= ptr_deref_860_load_2_req_0;
      reqL_unguarded(14) <= ptr_deref_819_load_1_req_0;
      reqL_unguarded(13) <= ptr_deref_807_load_2_req_0;
      reqL_unguarded(12) <= ptr_deref_807_load_3_req_0;
      reqL_unguarded(11) <= ptr_deref_976_load_0_req_0;
      reqL_unguarded(10) <= ptr_deref_976_load_1_req_0;
      reqL_unguarded(9) <= ptr_deref_976_load_2_req_0;
      reqL_unguarded(8) <= ptr_deref_976_load_3_req_0;
      reqL_unguarded(7) <= ptr_deref_1182_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_1182_load_1_req_0;
      reqL_unguarded(5) <= ptr_deref_1182_load_2_req_0;
      reqL_unguarded(4) <= ptr_deref_1182_load_3_req_0;
      reqL_unguarded(3) <= ptr_deref_1250_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1250_load_1_req_0;
      reqL_unguarded(1) <= ptr_deref_1250_load_2_req_0;
      reqL_unguarded(0) <= ptr_deref_1250_load_3_req_0;
      ptr_deref_819_load_3_ack_0 <= ackL_unguarded(23);
      ptr_deref_807_load_1_ack_0 <= ackL_unguarded(22);
      ptr_deref_819_load_2_ack_0 <= ackL_unguarded(21);
      ptr_deref_860_load_3_ack_0 <= ackL_unguarded(20);
      ptr_deref_860_load_1_ack_0 <= ackL_unguarded(19);
      ptr_deref_819_load_0_ack_0 <= ackL_unguarded(18);
      ptr_deref_807_load_0_ack_0 <= ackL_unguarded(17);
      ptr_deref_860_load_0_ack_0 <= ackL_unguarded(16);
      ptr_deref_860_load_2_ack_0 <= ackL_unguarded(15);
      ptr_deref_819_load_1_ack_0 <= ackL_unguarded(14);
      ptr_deref_807_load_2_ack_0 <= ackL_unguarded(13);
      ptr_deref_807_load_3_ack_0 <= ackL_unguarded(12);
      ptr_deref_976_load_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_976_load_1_ack_0 <= ackL_unguarded(10);
      ptr_deref_976_load_2_ack_0 <= ackL_unguarded(9);
      ptr_deref_976_load_3_ack_0 <= ackL_unguarded(8);
      ptr_deref_1182_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_1182_load_1_ack_0 <= ackL_unguarded(6);
      ptr_deref_1182_load_2_ack_0 <= ackL_unguarded(5);
      ptr_deref_1182_load_3_ack_0 <= ackL_unguarded(4);
      ptr_deref_1250_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1250_load_1_ack_0 <= ackL_unguarded(2);
      ptr_deref_1250_load_2_ack_0 <= ackL_unguarded(1);
      ptr_deref_1250_load_3_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(23) <= ptr_deref_819_load_3_req_1;
      reqR_unguarded(22) <= ptr_deref_807_load_1_req_1;
      reqR_unguarded(21) <= ptr_deref_819_load_2_req_1;
      reqR_unguarded(20) <= ptr_deref_860_load_3_req_1;
      reqR_unguarded(19) <= ptr_deref_860_load_1_req_1;
      reqR_unguarded(18) <= ptr_deref_819_load_0_req_1;
      reqR_unguarded(17) <= ptr_deref_807_load_0_req_1;
      reqR_unguarded(16) <= ptr_deref_860_load_0_req_1;
      reqR_unguarded(15) <= ptr_deref_860_load_2_req_1;
      reqR_unguarded(14) <= ptr_deref_819_load_1_req_1;
      reqR_unguarded(13) <= ptr_deref_807_load_2_req_1;
      reqR_unguarded(12) <= ptr_deref_807_load_3_req_1;
      reqR_unguarded(11) <= ptr_deref_976_load_0_req_1;
      reqR_unguarded(10) <= ptr_deref_976_load_1_req_1;
      reqR_unguarded(9) <= ptr_deref_976_load_2_req_1;
      reqR_unguarded(8) <= ptr_deref_976_load_3_req_1;
      reqR_unguarded(7) <= ptr_deref_1182_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_1182_load_1_req_1;
      reqR_unguarded(5) <= ptr_deref_1182_load_2_req_1;
      reqR_unguarded(4) <= ptr_deref_1182_load_3_req_1;
      reqR_unguarded(3) <= ptr_deref_1250_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1250_load_1_req_1;
      reqR_unguarded(1) <= ptr_deref_1250_load_2_req_1;
      reqR_unguarded(0) <= ptr_deref_1250_load_3_req_1;
      ptr_deref_819_load_3_ack_1 <= ackR_unguarded(23);
      ptr_deref_807_load_1_ack_1 <= ackR_unguarded(22);
      ptr_deref_819_load_2_ack_1 <= ackR_unguarded(21);
      ptr_deref_860_load_3_ack_1 <= ackR_unguarded(20);
      ptr_deref_860_load_1_ack_1 <= ackR_unguarded(19);
      ptr_deref_819_load_0_ack_1 <= ackR_unguarded(18);
      ptr_deref_807_load_0_ack_1 <= ackR_unguarded(17);
      ptr_deref_860_load_0_ack_1 <= ackR_unguarded(16);
      ptr_deref_860_load_2_ack_1 <= ackR_unguarded(15);
      ptr_deref_819_load_1_ack_1 <= ackR_unguarded(14);
      ptr_deref_807_load_2_ack_1 <= ackR_unguarded(13);
      ptr_deref_807_load_3_ack_1 <= ackR_unguarded(12);
      ptr_deref_976_load_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_976_load_1_ack_1 <= ackR_unguarded(10);
      ptr_deref_976_load_2_ack_1 <= ackR_unguarded(9);
      ptr_deref_976_load_3_ack_1 <= ackR_unguarded(8);
      ptr_deref_1182_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_1182_load_1_ack_1 <= ackR_unguarded(6);
      ptr_deref_1182_load_2_ack_1 <= ackR_unguarded(5);
      ptr_deref_1182_load_3_ack_1 <= ackR_unguarded(4);
      ptr_deref_1250_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1250_load_1_ack_1 <= ackR_unguarded(2);
      ptr_deref_1250_load_2_ack_1 <= ackR_unguarded(1);
      ptr_deref_1250_load_3_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_16: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_16", num_slots => 1) -- 
        port map (req => reqL_unregulated(16), -- 
          ack => ackL_unregulated(16),
          regulated_req => reqL(16),
          regulated_ack => ackL(16),
          release_req => reqR(16),
          release_ack => ackR(16),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_17: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_17", num_slots => 1) -- 
        port map (req => reqL_unregulated(17), -- 
          ack => ackL_unregulated(17),
          regulated_req => reqL(17),
          regulated_ack => ackL(17),
          release_req => reqR(17),
          release_ack => ackR(17),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_18: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_18", num_slots => 1) -- 
        port map (req => reqL_unregulated(18), -- 
          ack => ackL_unregulated(18),
          regulated_req => reqL(18),
          regulated_ack => ackL(18),
          release_req => reqR(18),
          release_ack => ackR(18),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_19: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_19", num_slots => 1) -- 
        port map (req => reqL_unregulated(19), -- 
          ack => ackL_unregulated(19),
          regulated_req => reqL(19),
          regulated_ack => ackL(19),
          release_req => reqR(19),
          release_ack => ackR(19),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_20: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_20", num_slots => 1) -- 
        port map (req => reqL_unregulated(20), -- 
          ack => ackL_unregulated(20),
          regulated_req => reqL(20),
          regulated_ack => ackL(20),
          release_req => reqR(20),
          release_ack => ackR(20),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_21: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_21", num_slots => 1) -- 
        port map (req => reqL_unregulated(21), -- 
          ack => ackL_unregulated(21),
          regulated_req => reqL(21),
          regulated_ack => ackL(21),
          release_req => reqR(21),
          release_ack => ackR(21),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_22: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_22", num_slots => 1) -- 
        port map (req => reqL_unregulated(22), -- 
          ack => ackL_unregulated(22),
          regulated_req => reqL(22),
          regulated_ack => ackL(22),
          release_req => reqR(22),
          release_ack => ackR(22),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_23: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_23", num_slots => 1) -- 
        port map (req => reqL_unregulated(23), -- 
          ack => ackL_unregulated(23),
          regulated_req => reqL(23),
          regulated_ack => ackL(23),
          release_req => reqR(23),
          release_ack => ackR(23),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 24, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_819_word_address_3 & ptr_deref_807_word_address_1 & ptr_deref_819_word_address_2 & ptr_deref_860_word_address_3 & ptr_deref_860_word_address_1 & ptr_deref_819_word_address_0 & ptr_deref_807_word_address_0 & ptr_deref_860_word_address_0 & ptr_deref_860_word_address_2 & ptr_deref_819_word_address_1 & ptr_deref_807_word_address_2 & ptr_deref_807_word_address_3 & ptr_deref_976_word_address_0 & ptr_deref_976_word_address_1 & ptr_deref_976_word_address_2 & ptr_deref_976_word_address_3 & ptr_deref_1182_word_address_0 & ptr_deref_1182_word_address_1 & ptr_deref_1182_word_address_2 & ptr_deref_1182_word_address_3 & ptr_deref_1250_word_address_0 & ptr_deref_1250_word_address_1 & ptr_deref_1250_word_address_2 & ptr_deref_1250_word_address_3;
      ptr_deref_819_data_3 <= data_out(191 downto 184);
      ptr_deref_807_data_1 <= data_out(183 downto 176);
      ptr_deref_819_data_2 <= data_out(175 downto 168);
      ptr_deref_860_data_3 <= data_out(167 downto 160);
      ptr_deref_860_data_1 <= data_out(159 downto 152);
      ptr_deref_819_data_0 <= data_out(151 downto 144);
      ptr_deref_807_data_0 <= data_out(143 downto 136);
      ptr_deref_860_data_0 <= data_out(135 downto 128);
      ptr_deref_860_data_2 <= data_out(127 downto 120);
      ptr_deref_819_data_1 <= data_out(119 downto 112);
      ptr_deref_807_data_2 <= data_out(111 downto 104);
      ptr_deref_807_data_3 <= data_out(103 downto 96);
      ptr_deref_976_data_0 <= data_out(95 downto 88);
      ptr_deref_976_data_1 <= data_out(87 downto 80);
      ptr_deref_976_data_2 <= data_out(79 downto 72);
      ptr_deref_976_data_3 <= data_out(71 downto 64);
      ptr_deref_1182_data_0 <= data_out(63 downto 56);
      ptr_deref_1182_data_1 <= data_out(55 downto 48);
      ptr_deref_1182_data_2 <= data_out(47 downto 40);
      ptr_deref_1182_data_3 <= data_out(39 downto 32);
      ptr_deref_1250_data_0 <= data_out(31 downto 24);
      ptr_deref_1250_data_1 <= data_out(23 downto 16);
      ptr_deref_1250_data_2 <= data_out(15 downto 8);
      ptr_deref_1250_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 9,
        num_reqs => 24,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(8 downto 0),
          mtag => memory_space_2_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 24,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_831_load_0 ptr_deref_843_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_831_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_843_load_0_req_0;
      ptr_deref_831_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_843_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_831_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_843_load_0_req_1;
      ptr_deref_831_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_843_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_831_word_address_0 & ptr_deref_843_word_address_0;
      ptr_deref_831_data_0 <= data_out(63 downto 32);
      ptr_deref_843_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared store operator group (0) : ptr_deref_1038_store_0 ptr_deref_1141_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1038_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1141_store_0_req_0;
      ptr_deref_1038_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1141_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1038_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1141_store_0_req_1;
      ptr_deref_1038_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1141_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1038_word_address_0 & ptr_deref_1141_word_address_0;
      data_in <= ptr_deref_1038_data_0 & ptr_deref_1141_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_starting_787_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_starting_787_inst_req_0;
      RPIPE_Block0_starting_787_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_starting_787_inst_req_1;
      RPIPE_Block0_starting_787_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_788 <= data_out(7 downto 0);
      Block0_starting_read_0_gI: SplitGuardInterface generic map(name => "Block0_starting_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block0_starting_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_starting_pipe_read_req(0),
          oack => Block0_starting_pipe_read_ack(0),
          odata => Block0_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_complete_1272_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_complete_1272_inst_req_0;
      WPIPE_Block0_complete_1272_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_complete_1272_inst_req_1;
      WPIPE_Block0_complete_1272_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_788;
      Block0_complete_write_0_gI: SplitGuardInterface generic map(name => "Block0_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_complete_pipe_write_req(0),
          oack => Block0_complete_pipe_write_ack(0),
          odata => Block0_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_A_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(17 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(43 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(8 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(37 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- declarations related to module zeropad3D_A
  component zeropad3D_A is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_A
  signal zeropad3D_A_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_A_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_A_start_req : std_logic;
  signal zeropad3D_A_start_ack : std_logic;
  signal zeropad3D_A_fin_req   : std_logic;
  signal zeropad3D_A_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_complete
  signal Block0_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_complete
  signal Block0_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_starting
  signal Block0_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_starting
  signal Block0_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 7),
      memory_space_3_lr_tag => memory_space_3_lr_tag(37 downto 19),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 32),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 2),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(17 downto 9),
      memory_space_2_lr_tag => memory_space_2_lr_tag(43 downto 22),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(15 downto 8),
      memory_space_2_lc_tag => memory_space_2_lc_tag(9 downto 5),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(8 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(7 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(21 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(6 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(0 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(7 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(17 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      Block0_complete_pipe_read_req => Block0_complete_pipe_read_req(0 downto 0),
      Block0_complete_pipe_read_ack => Block0_complete_pipe_read_ack(0 downto 0),
      Block0_complete_pipe_read_data => Block0_complete_pipe_read_data(7 downto 0),
      Block0_starting_pipe_write_req => Block0_starting_pipe_write_req(0 downto 0),
      Block0_starting_pipe_write_ack => Block0_starting_pipe_write_ack(0 downto 0),
      Block0_starting_pipe_write_data => Block0_starting_pipe_write_data(7 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  -- module zeropad3D_A
  zeropad3D_A_instance:zeropad3D_A-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_A_start_req,
      start_ack => zeropad3D_A_start_ack,
      fin_req => zeropad3D_A_fin_req,
      fin_ack => zeropad3D_A_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(8 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(21 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(7 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(4 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(6 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(0 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(17 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(7 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      Block0_starting_pipe_read_req => Block0_starting_pipe_read_req(0 downto 0),
      Block0_starting_pipe_read_ack => Block0_starting_pipe_read_ack(0 downto 0),
      Block0_starting_pipe_read_data => Block0_starting_pipe_read_data(7 downto 0),
      Block0_complete_pipe_write_req => Block0_complete_pipe_write_req(0 downto 0),
      Block0_complete_pipe_write_ack => Block0_complete_pipe_write_ack(0 downto 0),
      Block0_complete_pipe_write_data => Block0_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_A_tag_in,
      tag_out => zeropad3D_A_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_A_tag_in <= (others => '0');
  zeropad3D_A_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_A_start_req, start_ack => zeropad3D_A_start_ack,  fin_req => zeropad3D_A_fin_req,  fin_ack => zeropad3D_A_fin_ack);
  Block0_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_complete_pipe_read_req,
      read_ack => Block0_complete_pipe_read_ack,
      read_data => Block0_complete_pipe_read_data,
      write_req => Block0_complete_pipe_write_req,
      write_ack => Block0_complete_pipe_write_ack,
      write_data => Block0_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_starting_pipe_read_req,
      read_ack => Block0_starting_pipe_read_ack,
      read_data => Block0_starting_pipe_read_data,
      write_req => Block0_starting_pipe_write_req,
      write_ack => Block0_starting_pipe_write_ack,
      write_data => Block0_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 2,
      num_stores => 1,
      addr_width => 9,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 2,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
