-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_out_row_high_31_load_0_req_0 : boolean;
  signal LOAD_out_row_high_31_load_0_ack_0 : boolean;
  signal LOAD_out_row_high_31_load_0_req_1 : boolean;
  signal LOAD_out_row_high_31_load_0_ack_1 : boolean;
  signal type_cast_35_inst_req_0 : boolean;
  signal type_cast_35_inst_ack_0 : boolean;
  signal type_cast_35_inst_req_1 : boolean;
  signal type_cast_35_inst_ack_1 : boolean;
  signal LOAD_out_col_high_38_load_0_req_0 : boolean;
  signal LOAD_out_col_high_38_load_0_ack_0 : boolean;
  signal LOAD_out_col_high_38_load_0_req_1 : boolean;
  signal LOAD_out_col_high_38_load_0_ack_1 : boolean;
  signal type_cast_145_inst_req_0 : boolean;
  signal type_cast_145_inst_ack_0 : boolean;
  signal type_cast_145_inst_req_1 : boolean;
  signal type_cast_42_inst_req_0 : boolean;
  signal type_cast_42_inst_ack_0 : boolean;
  signal type_cast_42_inst_req_1 : boolean;
  signal type_cast_42_inst_ack_1 : boolean;
  signal LOAD_out_depth_high_45_load_0_req_0 : boolean;
  signal LOAD_out_depth_high_45_load_0_ack_0 : boolean;
  signal LOAD_out_depth_high_45_load_0_req_1 : boolean;
  signal LOAD_out_depth_high_45_load_0_ack_1 : boolean;
  signal type_cast_49_inst_req_0 : boolean;
  signal type_cast_49_inst_ack_0 : boolean;
  signal type_cast_49_inst_req_1 : boolean;
  signal type_cast_49_inst_ack_1 : boolean;
  signal if_stmt_74_branch_req_0 : boolean;
  signal if_stmt_74_branch_ack_1 : boolean;
  signal if_stmt_74_branch_ack_0 : boolean;
  signal type_cast_83_inst_req_0 : boolean;
  signal type_cast_83_inst_ack_0 : boolean;
  signal type_cast_83_inst_req_1 : boolean;
  signal type_cast_83_inst_ack_1 : boolean;
  signal type_cast_87_inst_req_0 : boolean;
  signal type_cast_87_inst_ack_0 : boolean;
  signal type_cast_87_inst_req_1 : boolean;
  signal type_cast_87_inst_ack_1 : boolean;
  signal type_cast_96_inst_req_0 : boolean;
  signal type_cast_96_inst_ack_0 : boolean;
  signal type_cast_96_inst_req_1 : boolean;
  signal type_cast_96_inst_ack_1 : boolean;
  signal array_obj_ref_136_index_offset_req_0 : boolean;
  signal array_obj_ref_136_index_offset_ack_0 : boolean;
  signal array_obj_ref_136_index_offset_req_1 : boolean;
  signal array_obj_ref_136_index_offset_ack_1 : boolean;
  signal addr_of_137_final_reg_req_0 : boolean;
  signal addr_of_137_final_reg_ack_0 : boolean;
  signal addr_of_137_final_reg_req_1 : boolean;
  signal addr_of_137_final_reg_ack_1 : boolean;
  signal ptr_deref_141_load_0_req_0 : boolean;
  signal ptr_deref_141_load_0_ack_0 : boolean;
  signal ptr_deref_141_load_0_req_1 : boolean;
  signal ptr_deref_141_load_0_ack_1 : boolean;
  signal type_cast_145_inst_ack_1 : boolean;
  signal type_cast_155_inst_req_0 : boolean;
  signal type_cast_155_inst_ack_0 : boolean;
  signal type_cast_155_inst_req_1 : boolean;
  signal type_cast_155_inst_ack_1 : boolean;
  signal type_cast_165_inst_req_0 : boolean;
  signal type_cast_165_inst_ack_0 : boolean;
  signal type_cast_165_inst_req_1 : boolean;
  signal type_cast_165_inst_ack_1 : boolean;
  signal type_cast_175_inst_req_0 : boolean;
  signal type_cast_175_inst_ack_0 : boolean;
  signal type_cast_175_inst_req_1 : boolean;
  signal type_cast_175_inst_ack_1 : boolean;
  signal type_cast_185_inst_req_0 : boolean;
  signal type_cast_185_inst_ack_0 : boolean;
  signal type_cast_185_inst_req_1 : boolean;
  signal type_cast_185_inst_ack_1 : boolean;
  signal type_cast_195_inst_req_0 : boolean;
  signal type_cast_195_inst_ack_0 : boolean;
  signal type_cast_195_inst_req_1 : boolean;
  signal type_cast_195_inst_ack_1 : boolean;
  signal type_cast_205_inst_req_0 : boolean;
  signal type_cast_205_inst_ack_0 : boolean;
  signal type_cast_205_inst_req_1 : boolean;
  signal type_cast_205_inst_ack_1 : boolean;
  signal type_cast_215_inst_req_0 : boolean;
  signal type_cast_215_inst_ack_0 : boolean;
  signal type_cast_215_inst_req_1 : boolean;
  signal type_cast_215_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_217_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_217_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_217_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_217_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_220_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_220_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_220_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_220_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_223_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_223_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_223_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_223_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_ack_1 : boolean;
  signal if_stmt_252_branch_req_0 : boolean;
  signal if_stmt_252_branch_ack_1 : boolean;
  signal if_stmt_252_branch_ack_0 : boolean;
  signal phi_stmt_124_req_0 : boolean;
  signal type_cast_130_inst_req_0 : boolean;
  signal type_cast_130_inst_ack_0 : boolean;
  signal type_cast_130_inst_req_1 : boolean;
  signal type_cast_130_inst_ack_1 : boolean;
  signal phi_stmt_124_req_1 : boolean;
  signal phi_stmt_124_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(77 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(77);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (50) 
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_29/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/branch_block_stmt_29__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_Update/cr
      -- 
    rr_72_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_72_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => LOAD_out_row_high_31_load_0_req_0); -- 
    cr_83_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_83_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => LOAD_out_row_high_31_load_0_req_1); -- 
    cr_102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => type_cast_35_inst_req_1); -- 
    rr_119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => LOAD_out_col_high_38_load_0_req_0); -- 
    cr_130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => LOAD_out_col_high_38_load_0_req_1); -- 
    cr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => type_cast_42_inst_req_1); -- 
    rr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => LOAD_out_depth_high_45_load_0_req_0); -- 
    cr_177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => LOAD_out_depth_high_45_load_0_req_1); -- 
    cr_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => type_cast_49_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Sample/word_access_start/word_0/ra
      -- 
    ra_73_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_row_high_31_load_0_ack_0, ack => sendOutput_CP_26_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (12) 
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/LOAD_out_row_high_31_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/LOAD_out_row_high_31_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/LOAD_out_row_high_31_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_row_high_31_Update/LOAD_out_row_high_31_Merge/merge_ack
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_Sample/rr
      -- 
    ca_84_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_row_high_31_load_0_ack_1, ack => sendOutput_CP_26_elements(2)); -- 
    rr_97_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_97_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(2), ack => type_cast_35_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_Sample/ra
      -- 
    ra_98_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_35_inst_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	13 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_35_Update/ca
      -- 
    ca_103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_35_inst_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Sample/word_access_start/word_0/ra
      -- 
    ra_120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_38_load_0_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/LOAD_out_col_high_38_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/LOAD_out_col_high_38_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/LOAD_out_col_high_38_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_col_high_38_Update/LOAD_out_col_high_38_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_Sample/rr
      -- 
    ca_131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_38_load_0_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    rr_144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(6), ack => type_cast_42_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_Sample/ra
      -- 
    ra_145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_42_inst_ack_0, ack => sendOutput_CP_26_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_42_Update/ca
      -- 
    ca_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_42_inst_ack_1, ack => sendOutput_CP_26_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Sample/word_access_start/word_0/ra
      -- 
    ra_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_45_load_0_ack_0, ack => sendOutput_CP_26_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/LOAD_out_depth_high_45_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/LOAD_out_depth_high_45_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/LOAD_out_depth_high_45_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/LOAD_out_depth_high_45_Update/LOAD_out_depth_high_45_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_Sample/rr
      -- 
    ca_178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_45_load_0_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    rr_191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_49_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_Sample/ra
      -- 
    ra_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_49_inst_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/type_cast_49_Update/ca
      -- 
    ca_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_49_inst_ack_1, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  branch  join  transition  place  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: 	4 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (10) 
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73__exit__
      -- CP-element group 13: 	 branch_block_stmt_29/if_stmt_74__entry__
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_32_to_assign_stmt_73/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/if_stmt_74_dead_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/if_stmt_74_eval_test/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/if_stmt_74_eval_test/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/if_stmt_74_eval_test/branch_req
      -- CP-element group 13: 	 branch_block_stmt_29/R_cmp81_75_place
      -- CP-element group 13: 	 branch_block_stmt_29/if_stmt_74_if_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/if_stmt_74_else_link/$entry
      -- 
    branch_req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(13), ack => if_stmt_74_branch_req_0); -- 
    sendOutput_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(12) & sendOutput_CP_26_elements(4) & sendOutput_CP_26_elements(8);
      gj_sendOutput_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  transition  place  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	77 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_29/if_stmt_74_if_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_29/if_stmt_74_if_link/if_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_29/entry_forx_xend
      -- CP-element group 14: 	 branch_block_stmt_29/entry_forx_xend_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_29/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_74_branch_ack_1, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15:  members (30) 
      -- CP-element group 15: 	 branch_block_stmt_29/merge_stmt_80__exit__
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121__entry__
      -- CP-element group 15: 	 branch_block_stmt_29/if_stmt_74_else_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/if_stmt_74_else_link/else_choice_transition
      -- CP-element group 15: 	 branch_block_stmt_29/entry_bbx_xnph
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_update_start_
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_update_start_
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_update_start_
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_29/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/merge_stmt_80_PhiReqMerge
      -- CP-element group 15: 	 branch_block_stmt_29/merge_stmt_80_PhiAck/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/merge_stmt_80_PhiAck/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/merge_stmt_80_PhiAck/dummy
      -- 
    else_choice_transition_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_74_branch_ack_0, ack => sendOutput_CP_26_elements(15)); -- 
    rr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => type_cast_83_inst_req_0); -- 
    cr_232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => type_cast_83_inst_req_1); -- 
    rr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => type_cast_87_inst_req_0); -- 
    cr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => type_cast_87_inst_req_1); -- 
    rr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => type_cast_96_inst_req_0); -- 
    cr_260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => type_cast_96_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_Sample/ra
      -- 
    ra_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_0, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	22 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_83_Update/ca
      -- 
    ca_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_1, ack => sendOutput_CP_26_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_Sample/ra
      -- 
    ra_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_87_inst_ack_0, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_87_Update/ca
      -- 
    ca_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_87_inst_ack_1, ack => sendOutput_CP_26_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_Sample/ra
      -- 
    ra_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_96_inst_ack_0, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/type_cast_96_Update/ca
      -- 
    ca_261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_96_inst_ack_1, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  join  transition  place  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	17 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	71 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121__exit__
      -- CP-element group 22: 	 branch_block_stmt_29/bbx_xnph_forx_xbody
      -- CP-element group 22: 	 branch_block_stmt_29/assign_stmt_84_to_assign_stmt_121/$exit
      -- CP-element group 22: 	 branch_block_stmt_29/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 22: 	 branch_block_stmt_29/bbx_xnph_forx_xbody_PhiReq/phi_stmt_124/$entry
      -- CP-element group 22: 	 branch_block_stmt_29/bbx_xnph_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/$entry
      -- 
    sendOutput_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(17) & sendOutput_CP_26_elements(19) & sendOutput_CP_26_elements(21);
      gj_sendOutput_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	76 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	68 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_sample_complete
      -- CP-element group 23: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_Sample/ack
      -- 
    ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_136_index_offset_ack_0, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	76 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (11) 
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_root_address_calculated
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_offset_calculated
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_Update/ack
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_base_plus_offset/$entry
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_base_plus_offset/$exit
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_base_plus_offset/sum_rename_req
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_base_plus_offset/sum_rename_ack
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_request/$entry
      -- CP-element group 24: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_request/req
      -- 
    ack_295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_136_index_offset_ack_1, ack => sendOutput_CP_26_elements(24)); -- 
    req_304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(24), ack => addr_of_137_final_reg_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_request/$exit
      -- CP-element group 25: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_request/ack
      -- 
    ack_305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_137_final_reg_ack_0, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	76 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (24) 
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_complete/ack
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_word_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_root_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_address_resized
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_addr_resize/$entry
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_addr_resize/$exit
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_addr_resize/base_resize_req
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_addr_resize/base_resize_ack
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_plus_offset/$entry
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_plus_offset/$exit
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_base_plus_offset/sum_rename_ack
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_word_addrgen/$entry
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_word_addrgen/$exit
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_word_addrgen/root_register_req
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_word_addrgen/root_register_ack
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Sample/word_access_start/$entry
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Sample/word_access_start/word_0/$entry
      -- CP-element group 26: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Sample/word_access_start/word_0/rr
      -- 
    ack_310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_137_final_reg_ack_1, ack => sendOutput_CP_26_elements(26)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(26), ack => ptr_deref_141_load_0_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Sample/word_access_start/word_0/ra
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_141_load_0_ack_0, ack => sendOutput_CP_26_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	76 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	31 
    -- CP-element group 28: 	33 
    -- CP-element group 28: 	35 
    -- CP-element group 28: 	37 
    -- CP-element group 28: 	39 
    -- CP-element group 28: 	41 
    -- CP-element group 28: 	43 
    -- CP-element group 28:  members (33) 
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/ptr_deref_141_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/ptr_deref_141_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/ptr_deref_141_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/ptr_deref_141_Merge/merge_ack
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_Sample/rr
      -- 
    ca_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_141_load_0_ack_1, ack => sendOutput_CP_26_elements(28)); -- 
    rr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(28), ack => type_cast_145_inst_req_0); -- 
    rr_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(28), ack => type_cast_155_inst_req_0); -- 
    rr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(28), ack => type_cast_165_inst_req_0); -- 
    rr_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(28), ack => type_cast_175_inst_req_0); -- 
    rr_424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(28), ack => type_cast_185_inst_req_0); -- 
    rr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(28), ack => type_cast_195_inst_req_0); -- 
    rr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(28), ack => type_cast_205_inst_req_0); -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(28), ack => type_cast_215_inst_req_0); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_Sample/ra
      -- 
    ra_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_0, ack => sendOutput_CP_26_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	76 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	65 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_Update/ca
      -- 
    ca_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_1, ack => sendOutput_CP_26_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	28 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_Sample/ra
      -- 
    ra_383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_0, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	76 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	62 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_Update/ca
      -- 
    ca_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_1, ack => sendOutput_CP_26_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	28 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_Sample/ra
      -- 
    ra_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_165_inst_ack_0, ack => sendOutput_CP_26_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	76 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	59 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_Update/ca
      -- 
    ca_402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_165_inst_ack_1, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	28 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_Sample/ra
      -- 
    ra_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_175_inst_ack_0, ack => sendOutput_CP_26_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	76 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	56 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_Update/ca
      -- 
    ca_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_175_inst_ack_1, ack => sendOutput_CP_26_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	28 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_Sample/ra
      -- 
    ra_425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_0, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	76 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	53 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_Update/ca
      -- 
    ca_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_1, ack => sendOutput_CP_26_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	28 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_Sample/ra
      -- 
    ra_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	76 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	50 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_Update/ca
      -- 
    ca_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	28 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_Sample/ra
      -- 
    ra_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_0, ack => sendOutput_CP_26_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	76 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	47 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_Update/ca
      -- 
    ca_458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_1, ack => sendOutput_CP_26_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	28 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_0, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	76 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_Sample/req
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_1, ack => sendOutput_CP_26_elements(44)); -- 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_217_inst_req_0); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_update_start_
      -- CP-element group 45: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_Update/req
      -- 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_217_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_217_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_217_Update/ack
      -- 
    ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_217_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	42 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_Sample/req
      -- 
    req_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_220_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(42) & sendOutput_CP_26_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_update_start_
      -- CP-element group 48: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_Update/req
      -- 
    ack_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_220_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_220_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_220_Update/ack
      -- 
    ack_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_220_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	40 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_Sample/req
      -- 
    req_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => WPIPE_zeropad_output_pipe_223_inst_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(40) & sendOutput_CP_26_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_update_start_
      -- CP-element group 51: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_Update/req
      -- 
    ack_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_223_inst_ack_0, ack => sendOutput_CP_26_elements(51)); -- 
    req_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(51), ack => WPIPE_zeropad_output_pipe_223_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_223_Update/ack
      -- 
    ack_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_223_inst_ack_1, ack => sendOutput_CP_26_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	38 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_Sample/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => WPIPE_zeropad_output_pipe_226_inst_req_0); -- 
    sendOutput_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(38) & sendOutput_CP_26_elements(52);
      gj_sendOutput_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_update_start_
      -- CP-element group 54: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_Update/req
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_226_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(54), ack => WPIPE_zeropad_output_pipe_226_inst_req_1); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_226_Update/ack
      -- 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_226_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_Sample/req
      -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => WPIPE_zeropad_output_pipe_229_inst_req_0); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(36) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_update_start_
      -- CP-element group 57: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_Update/req
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_229_inst_ack_0, ack => sendOutput_CP_26_elements(57)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(57), ack => WPIPE_zeropad_output_pipe_229_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_229_Update/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_229_inst_ack_1, ack => sendOutput_CP_26_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	34 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_Sample/req
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(59), ack => WPIPE_zeropad_output_pipe_232_inst_req_0); -- 
    sendOutput_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(34) & sendOutput_CP_26_elements(58);
      gj_sendOutput_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_update_start_
      -- CP-element group 60: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_Update/req
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_232_inst_ack_0, ack => sendOutput_CP_26_elements(60)); -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(60), ack => WPIPE_zeropad_output_pipe_232_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_232_Update/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_232_inst_ack_1, ack => sendOutput_CP_26_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	32 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_Sample/req
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(62), ack => WPIPE_zeropad_output_pipe_235_inst_req_0); -- 
    sendOutput_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(32) & sendOutput_CP_26_elements(61);
      gj_sendOutput_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_update_start_
      -- CP-element group 63: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_Update/req
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_235_inst_ack_0, ack => sendOutput_CP_26_elements(63)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(63), ack => WPIPE_zeropad_output_pipe_235_inst_req_1); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_235_Update/ack
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_235_inst_ack_1, ack => sendOutput_CP_26_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	30 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_Sample/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(65), ack => WPIPE_zeropad_output_pipe_238_inst_req_0); -- 
    sendOutput_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(30) & sendOutput_CP_26_elements(64);
      gj_sendOutput_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_update_start_
      -- CP-element group 66: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_Update/req
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_238_inst_ack_0, ack => sendOutput_CP_26_elements(66)); -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(66), ack => WPIPE_zeropad_output_pipe_238_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/WPIPE_zeropad_output_pipe_238_Update/ack
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_238_inst_ack_1, ack => sendOutput_CP_26_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	23 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251__exit__
      -- CP-element group 68: 	 branch_block_stmt_29/if_stmt_252__entry__
      -- CP-element group 68: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/$exit
      -- CP-element group 68: 	 branch_block_stmt_29/if_stmt_252_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_29/if_stmt_252_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_29/if_stmt_252_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_29/if_stmt_252_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_29/R_exitcond11_253_place
      -- CP-element group 68: 	 branch_block_stmt_29/if_stmt_252_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_29/if_stmt_252_else_link/$entry
      -- 
    branch_req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(68), ack => if_stmt_252_branch_req_0); -- 
    sendOutput_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(23) & sendOutput_CP_26_elements(67);
      gj_sendOutput_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  transition  place  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	77 
    -- CP-element group 69:  members (13) 
      -- CP-element group 69: 	 branch_block_stmt_29/merge_stmt_258__exit__
      -- CP-element group 69: 	 branch_block_stmt_29/forx_xendx_xloopexit_forx_xend
      -- CP-element group 69: 	 branch_block_stmt_29/if_stmt_252_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_29/if_stmt_252_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_29/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 69: 	 branch_block_stmt_29/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_29/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_29/merge_stmt_258_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_29/merge_stmt_258_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_29/merge_stmt_258_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_29/merge_stmt_258_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_29/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_29/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_252_branch_ack_1, ack => sendOutput_CP_26_elements(69)); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	73 
    -- CP-element group 70:  members (12) 
      -- CP-element group 70: 	 branch_block_stmt_29/if_stmt_252_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_29/if_stmt_252_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/$entry
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/$entry
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/Update/cr
      -- 
    else_choice_transition_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_252_branch_ack_0, ack => sendOutput_CP_26_elements(70)); -- 
    rr_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(70), ack => type_cast_130_inst_req_0); -- 
    cr_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(70), ack => type_cast_130_inst_req_1); -- 
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	22 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_29/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_29/bbx_xnph_forx_xbody_PhiReq/phi_stmt_124/$exit
      -- CP-element group 71: 	 branch_block_stmt_29/bbx_xnph_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_29/bbx_xnph_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_128_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_29/bbx_xnph_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_req
      -- 
    phi_stmt_124_req_626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_124_req_626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(71), ack => phi_stmt_124_req_0); -- 
    -- Element group sendOutput_CP_26_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(22), ack => sendOutput_CP_26_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/Sample/ra
      -- 
    ra_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_130_inst_ack_0, ack => sendOutput_CP_26_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	70 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/Update/ca
      -- 
    ca_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_130_inst_ack_1, ack => sendOutput_CP_26_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/$exit
      -- CP-element group 74: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/$exit
      -- CP-element group 74: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_sources/type_cast_130/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_29/forx_xbody_forx_xbody_PhiReq/phi_stmt_124/phi_stmt_124_req
      -- 
    phi_stmt_124_req_652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_124_req_652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(74), ack => phi_stmt_124_req_1); -- 
    sendOutput_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(72) & sendOutput_CP_26_elements(73);
      gj_sendOutput_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  transition  place  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_29/merge_stmt_123_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_29/merge_stmt_123_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(75) <= OrReduce(sendOutput_CP_26_elements(71) & sendOutput_CP_26_elements(74));
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	23 
    -- CP-element group 76: 	24 
    -- CP-element group 76: 	26 
    -- CP-element group 76: 	28 
    -- CP-element group 76: 	30 
    -- CP-element group 76: 	32 
    -- CP-element group 76: 	34 
    -- CP-element group 76: 	36 
    -- CP-element group 76: 	38 
    -- CP-element group 76: 	40 
    -- CP-element group 76: 	42 
    -- CP-element group 76: 	44 
    -- CP-element group 76:  members (53) 
      -- CP-element group 76: 	 branch_block_stmt_29/merge_stmt_123__exit__
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251__entry__
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_145_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_resized_1
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_scaled_1
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_computed_1
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_resize_1/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_resize_1/$exit
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_resize_1/index_resize_req
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_resize_1/index_resize_ack
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_scale_1/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_scale_1/$exit
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_scale_1/scale_rename_req
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_index_scale_1/scale_rename_ack
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_update_start
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_Sample/req
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/array_obj_ref_136_final_index_sum_regn_Update/req
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_complete/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/addr_of_137_complete/req
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/word_access_complete/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/word_access_complete/word_0/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/ptr_deref_141_Update/word_access_complete/word_0/cr
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_155_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_165_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_175_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_185_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_195_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_205_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_update_start_
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_29/assign_stmt_138_to_assign_stmt_251/type_cast_215_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_29/merge_stmt_123_PhiAck/$exit
      -- CP-element group 76: 	 branch_block_stmt_29/merge_stmt_123_PhiAck/phi_stmt_124_ack
      -- 
    phi_stmt_124_ack_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_124_ack_0, ack => sendOutput_CP_26_elements(76)); -- 
    cr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => type_cast_145_inst_req_1); -- 
    req_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => array_obj_ref_136_index_offset_req_0); -- 
    req_294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => array_obj_ref_136_index_offset_req_1); -- 
    req_309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => addr_of_137_final_reg_req_1); -- 
    cr_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => ptr_deref_141_load_0_req_1); -- 
    cr_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => type_cast_155_inst_req_1); -- 
    cr_401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => type_cast_165_inst_req_1); -- 
    cr_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => type_cast_175_inst_req_1); -- 
    cr_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => type_cast_185_inst_req_1); -- 
    cr_443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => type_cast_195_inst_req_1); -- 
    cr_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => type_cast_205_inst_req_1); -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(76), ack => type_cast_215_inst_req_1); -- 
    -- CP-element group 77:  merge  transition  place  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	14 
    -- CP-element group 77: 	69 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (16) 
      -- CP-element group 77: 	 $exit
      -- CP-element group 77: 	 branch_block_stmt_29/$exit
      -- CP-element group 77: 	 branch_block_stmt_29/branch_block_stmt_29__exit__
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_260__exit__
      -- CP-element group 77: 	 branch_block_stmt_29/return__
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_262__exit__
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_260_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_260_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_260_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_260_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_29/return___PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_29/return___PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_262_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_262_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_262_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_29/merge_stmt_262_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(77) <= OrReduce(sendOutput_CP_26_elements(14) & sendOutput_CP_26_elements(69));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_out_col_high_38_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_38_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_45_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_45_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_row_high_31_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_row_high_31_word_address_0 : std_logic_vector(0 downto 0);
    signal R_indvar_135_resized : std_logic_vector(13 downto 0);
    signal R_indvar_135_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_136_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_136_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_136_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_136_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_136_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_136_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_138 : std_logic_vector(31 downto 0);
    signal cmp81_73 : std_logic_vector(0 downto 0);
    signal conv17_146 : std_logic_vector(7 downto 0);
    signal conv23_156 : std_logic_vector(7 downto 0);
    signal conv29_166 : std_logic_vector(7 downto 0);
    signal conv2_43 : std_logic_vector(63 downto 0);
    signal conv35_176 : std_logic_vector(7 downto 0);
    signal conv41_186 : std_logic_vector(7 downto 0);
    signal conv47_196 : std_logic_vector(7 downto 0);
    signal conv4_50 : std_logic_vector(63 downto 0);
    signal conv53_206 : std_logic_vector(7 downto 0);
    signal conv59_216 : std_logic_vector(7 downto 0);
    signal conv_36 : std_logic_vector(63 downto 0);
    signal exitcond11_251 : std_logic_vector(0 downto 0);
    signal indvar_124 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_246 : std_logic_vector(63 downto 0);
    signal mul5_60 : std_logic_vector(63 downto 0);
    signal mul_55 : std_logic_vector(63 downto 0);
    signal ptr_deref_141_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_141_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_141_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_141_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_141_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr20_152 : std_logic_vector(63 downto 0);
    signal shr26_162 : std_logic_vector(63 downto 0);
    signal shr32_172 : std_logic_vector(63 downto 0);
    signal shr38_182 : std_logic_vector(63 downto 0);
    signal shr44_192 : std_logic_vector(63 downto 0);
    signal shr50_202 : std_logic_vector(63 downto 0);
    signal shr56_212 : std_logic_vector(63 downto 0);
    signal shr80x_xmask_66 : std_logic_vector(63 downto 0);
    signal tmp14_142 : std_logic_vector(63 downto 0);
    signal tmp1_39 : std_logic_vector(7 downto 0);
    signal tmp2_84 : std_logic_vector(63 downto 0);
    signal tmp3_46 : std_logic_vector(7 downto 0);
    signal tmp4_88 : std_logic_vector(63 downto 0);
    signal tmp5_93 : std_logic_vector(63 downto 0);
    signal tmp6_97 : std_logic_vector(63 downto 0);
    signal tmp7_102 : std_logic_vector(63 downto 0);
    signal tmp8_108 : std_logic_vector(63 downto 0);
    signal tmp9_114 : std_logic_vector(0 downto 0);
    signal tmp_32 : std_logic_vector(7 downto 0);
    signal type_cast_106_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_112_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_119_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_128_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_130_wire : std_logic_vector(63 downto 0);
    signal type_cast_150_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_160_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_170_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_180_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_190_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_200_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_210_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_244_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_64_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_70_wire_constant : std_logic_vector(63 downto 0);
    signal umax10_121 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    LOAD_out_col_high_38_word_address_0 <= "0";
    LOAD_out_depth_high_45_word_address_0 <= "0";
    LOAD_out_row_high_31_word_address_0 <= "0";
    array_obj_ref_136_constant_part_of_offset <= "00000000000000";
    array_obj_ref_136_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_136_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_136_resized_base_address <= "00000000000000";
    ptr_deref_141_word_offset_0 <= "00000000000000";
    type_cast_106_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_119_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_128_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_150_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_160_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_170_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_180_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_190_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_200_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_210_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_244_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_64_wire_constant <= "0000000000000000000000000000000000000000111111111111111111111100";
    type_cast_70_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_124: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_128_wire_constant & type_cast_130_wire;
      req <= phi_stmt_124_req_0 & phi_stmt_124_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_124",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_124_ack_0,
          idata => idata,
          odata => indvar_124,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_124
    -- flow-through select operator MUX_120_inst
    umax10_121 <= tmp8_108 when (tmp9_114(0) /=  '0') else type_cast_119_wire_constant;
    addr_of_137_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_137_final_reg_req_0;
      addr_of_137_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_137_final_reg_req_1;
      addr_of_137_final_reg_ack_1<= rack(0);
      addr_of_137_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_137_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_136_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_138,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_130_inst_req_0;
      type_cast_130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_130_inst_req_1;
      type_cast_130_inst_ack_1<= rack(0);
      type_cast_130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_130_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_145_inst_req_0;
      type_cast_145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_145_inst_req_1;
      type_cast_145_inst_ack_1<= rack(0);
      type_cast_145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_155_inst_req_0;
      type_cast_155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_155_inst_req_1;
      type_cast_155_inst_ack_1<= rack(0);
      type_cast_155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr20_152,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_156,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_165_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_165_inst_req_0;
      type_cast_165_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_165_inst_req_1;
      type_cast_165_inst_ack_1<= rack(0);
      type_cast_165_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_165_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr26_162,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_166,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_175_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_175_inst_req_0;
      type_cast_175_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_175_inst_req_1;
      type_cast_175_inst_ack_1<= rack(0);
      type_cast_175_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_175_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr32_172,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_176,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_185_inst_req_0;
      type_cast_185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_185_inst_req_1;
      type_cast_185_inst_ack_1<= rack(0);
      type_cast_185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr38_182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_186,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_195_inst_req_0;
      type_cast_195_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_195_inst_req_1;
      type_cast_195_inst_ack_1<= rack(0);
      type_cast_195_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_195_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr44_192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_205_inst_req_0;
      type_cast_205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_205_inst_req_1;
      type_cast_205_inst_ack_1<= rack(0);
      type_cast_205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr50_202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_215_inst_req_0;
      type_cast_215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_215_inst_req_1;
      type_cast_215_inst_ack_1<= rack(0);
      type_cast_215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr56_212,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_35_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_35_inst_req_0;
      type_cast_35_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_35_inst_req_1;
      type_cast_35_inst_ack_1<= rack(0);
      type_cast_35_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_35_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_32,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_36,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_42_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_42_inst_req_0;
      type_cast_42_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_42_inst_req_1;
      type_cast_42_inst_ack_1<= rack(0);
      type_cast_42_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_42_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_39,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_43,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_49_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_49_inst_req_0;
      type_cast_49_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_49_inst_req_1;
      type_cast_49_inst_ack_1<= rack(0);
      type_cast_49_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_49_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_46,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_50,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_83_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_83_inst_req_0;
      type_cast_83_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_83_inst_req_1;
      type_cast_83_inst_ack_1<= rack(0);
      type_cast_83_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_83_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_39,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp2_84,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_87_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_87_inst_req_0;
      type_cast_87_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_87_inst_req_1;
      type_cast_87_inst_ack_1<= rack(0);
      type_cast_87_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_87_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_32,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp4_88,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_96_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_96_inst_req_0;
      type_cast_96_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_96_inst_req_1;
      type_cast_96_inst_ack_1<= rack(0);
      type_cast_96_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_96_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_46,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_97,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_out_col_high_38_gather_scatter
    process(LOAD_out_col_high_38_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_38_data_0;
      ov(7 downto 0) := iv;
      tmp1_39 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_45_gather_scatter
    process(LOAD_out_depth_high_45_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_45_data_0;
      ov(7 downto 0) := iv;
      tmp3_46 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_row_high_31_gather_scatter
    process(LOAD_out_row_high_31_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_row_high_31_data_0;
      ov(7 downto 0) := iv;
      tmp_32 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_136_index_1_rename
    process(R_indvar_135_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_135_resized;
      ov(13 downto 0) := iv;
      R_indvar_135_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_136_index_1_resize
    process(indvar_124) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_124;
      ov := iv(13 downto 0);
      R_indvar_135_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_136_root_address_inst
    process(array_obj_ref_136_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_136_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_136_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_141_addr_0
    process(ptr_deref_141_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_141_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_141_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_141_base_resize
    process(arrayidx_138) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_138;
      ov := iv(13 downto 0);
      ptr_deref_141_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_141_gather_scatter
    process(ptr_deref_141_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_141_data_0;
      ov(63 downto 0) := iv;
      tmp14_142 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_141_root_address_inst
    process(ptr_deref_141_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_141_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_141_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_252_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond11_251;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_252_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_252_branch_req_0,
          ack0 => if_stmt_252_branch_ack_0,
          ack1 => if_stmt_252_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_74_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp81_73;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_74_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_74_branch_req_0,
          ack0 => if_stmt_74_branch_ack_0,
          ack1 => if_stmt_74_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_245_inst
    process(indvar_124) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_124, type_cast_244_wire_constant, tmp_var);
      indvarx_xnext_246 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_65_inst
    process(mul5_60) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul5_60, type_cast_64_wire_constant, tmp_var);
      shr80x_xmask_66 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_250_inst
    process(indvarx_xnext_246, umax10_121) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_246, umax10_121, tmp_var);
      exitcond11_251 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_71_inst
    process(shr80x_xmask_66) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr80x_xmask_66, type_cast_70_wire_constant, tmp_var);
      cmp81_73 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_107_inst
    process(tmp7_102) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp7_102, type_cast_106_wire_constant, tmp_var);
      tmp8_108 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_151_inst
    process(tmp14_142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_142, type_cast_150_wire_constant, tmp_var);
      shr20_152 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_161_inst
    process(tmp14_142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_142, type_cast_160_wire_constant, tmp_var);
      shr26_162 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_171_inst
    process(tmp14_142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_142, type_cast_170_wire_constant, tmp_var);
      shr32_172 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_181_inst
    process(tmp14_142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_142, type_cast_180_wire_constant, tmp_var);
      shr38_182 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_191_inst
    process(tmp14_142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_142, type_cast_190_wire_constant, tmp_var);
      shr44_192 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_201_inst
    process(tmp14_142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_142, type_cast_200_wire_constant, tmp_var);
      shr50_202 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_211_inst
    process(tmp14_142) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_142, type_cast_210_wire_constant, tmp_var);
      shr56_212 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_101_inst
    process(tmp5_93, tmp6_97) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp5_93, tmp6_97, tmp_var);
      tmp7_102 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_54_inst
    process(conv2_43, conv_36) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv2_43, conv_36, tmp_var);
      mul_55 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_59_inst
    process(mul_55, conv4_50) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_55, conv4_50, tmp_var);
      mul5_60 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_92_inst
    process(tmp2_84, tmp4_88) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_84, tmp4_88, tmp_var);
      tmp5_93 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_113_inst
    process(tmp8_108) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp8_108, type_cast_112_wire_constant, tmp_var);
      tmp9_114 <= tmp_var; --
    end process;
    -- shared split operator group (17) : array_obj_ref_136_index_offset 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_135_scaled;
      array_obj_ref_136_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_136_index_offset_req_0;
      array_obj_ref_136_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_136_index_offset_req_1;
      array_obj_ref_136_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared load operator group (0) : LOAD_out_col_high_38_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_out_col_high_38_load_0_req_0;
      LOAD_out_col_high_38_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_out_col_high_38_load_0_req_1;
      LOAD_out_col_high_38_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_out_col_high_38_word_address_0;
      LOAD_out_col_high_38_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(7 downto 0),
          mtag => memory_space_6_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : LOAD_out_depth_high_45_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_out_depth_high_45_load_0_req_0;
      LOAD_out_depth_high_45_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_out_depth_high_45_load_0_req_1;
      LOAD_out_depth_high_45_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_out_depth_high_45_word_address_0;
      LOAD_out_depth_high_45_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : LOAD_out_row_high_31_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_out_row_high_31_load_0_req_0;
      LOAD_out_row_high_31_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_out_row_high_31_load_0_req_1;
      LOAD_out_row_high_31_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_out_row_high_31_word_address_0;
      LOAD_out_row_high_31_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(7 downto 0),
          mtag => memory_space_8_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_141_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_141_load_0_req_0;
      ptr_deref_141_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_141_load_0_req_1;
      ptr_deref_141_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_141_word_address_0;
      ptr_deref_141_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 14,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_217_inst WPIPE_zeropad_output_pipe_220_inst WPIPE_zeropad_output_pipe_223_inst WPIPE_zeropad_output_pipe_226_inst WPIPE_zeropad_output_pipe_229_inst WPIPE_zeropad_output_pipe_232_inst WPIPE_zeropad_output_pipe_235_inst WPIPE_zeropad_output_pipe_238_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_217_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_220_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_223_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_226_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_229_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_232_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_235_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_238_inst_req_0;
      WPIPE_zeropad_output_pipe_217_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_220_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_223_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_226_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_229_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_232_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_235_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_238_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_217_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_220_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_223_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_226_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_229_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_232_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_235_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_238_inst_req_1;
      WPIPE_zeropad_output_pipe_217_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_220_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_223_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_226_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_229_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_232_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_235_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_238_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv59_216 & conv53_206 & conv47_196 & conv41_186 & conv35_176 & conv29_166 & conv23_156 & conv17_146;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_10_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_10_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_9_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_9_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_10_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_10_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_689_start: Boolean;
  signal testConfigure_CP_689_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_zeropad_input_pipe_321_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_321_inst_ack_1 : boolean;
  signal ptr_deref_311_store_0_ack_1 : boolean;
  signal STORE_col_high_323_store_0_req_0 : boolean;
  signal type_cast_590_inst_ack_0 : boolean;
  signal STORE_col_high_323_store_0_ack_0 : boolean;
  signal type_cast_623_inst_ack_0 : boolean;
  signal phi_stmt_449_req_0 : boolean;
  signal ptr_deref_598_store_0_ack_1 : boolean;
  signal type_cast_590_inst_ack_1 : boolean;
  signal type_cast_590_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_281_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_321_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_281_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_298_inst_ack_1 : boolean;
  signal type_cast_285_inst_ack_1 : boolean;
  signal STORE_row_high_317_store_0_ack_1 : boolean;
  signal type_cast_285_inst_req_1 : boolean;
  signal STORE_row_high_317_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_298_inst_req_1 : boolean;
  signal type_cast_482_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_298_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_298_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_315_inst_ack_1 : boolean;
  signal phi_stmt_449_req_1 : boolean;
  signal type_cast_285_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_315_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_281_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_281_inst_req_0 : boolean;
  signal type_cast_285_inst_req_0 : boolean;
  signal type_cast_500_inst_ack_0 : boolean;
  signal type_cast_518_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_550_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_315_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_315_inst_req_0 : boolean;
  signal type_cast_455_inst_ack_1 : boolean;
  signal ptr_deref_276_store_0_ack_1 : boolean;
  signal type_cast_482_inst_ack_0 : boolean;
  signal type_cast_482_inst_req_1 : boolean;
  signal ptr_deref_276_store_0_req_1 : boolean;
  signal ptr_deref_294_store_0_ack_1 : boolean;
  signal ptr_deref_294_store_0_req_1 : boolean;
  signal STORE_row_high_317_store_0_ack_0 : boolean;
  signal STORE_row_high_317_store_0_req_0 : boolean;
  signal ptr_deref_311_store_0_req_1 : boolean;
  signal ptr_deref_294_store_0_ack_0 : boolean;
  signal ptr_deref_276_store_0_ack_0 : boolean;
  signal ptr_deref_294_store_0_req_0 : boolean;
  signal type_cast_518_inst_req_0 : boolean;
  signal ptr_deref_276_store_0_req_0 : boolean;
  signal type_cast_623_inst_req_1 : boolean;
  signal type_cast_518_inst_ack_0 : boolean;
  signal type_cast_518_inst_req_1 : boolean;
  signal type_cast_623_inst_ack_1 : boolean;
  signal type_cast_302_inst_ack_1 : boolean;
  signal type_cast_302_inst_req_1 : boolean;
  signal type_cast_302_inst_ack_0 : boolean;
  signal type_cast_302_inst_req_0 : boolean;
  signal ptr_deref_311_store_0_ack_0 : boolean;
  signal ptr_deref_311_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_321_inst_req_0 : boolean;
  signal type_cast_455_inst_req_1 : boolean;
  signal type_cast_500_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_550_inst_ack_1 : boolean;
  signal type_cast_482_inst_ack_1 : boolean;
  signal if_stmt_612_branch_req_0 : boolean;
  signal type_cast_500_inst_req_1 : boolean;
  signal type_cast_500_inst_ack_1 : boolean;
  signal if_stmt_612_branch_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_532_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_532_inst_ack_0 : boolean;
  signal ptr_deref_598_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_532_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_532_inst_ack_1 : boolean;
  signal ptr_deref_598_store_0_ack_0 : boolean;
  signal if_stmt_612_branch_ack_0 : boolean;
  signal phi_stmt_449_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_496_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_496_inst_ack_0 : boolean;
  signal type_cast_536_inst_req_0 : boolean;
  signal type_cast_455_inst_req_0 : boolean;
  signal ptr_deref_598_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_496_inst_req_1 : boolean;
  signal type_cast_536_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_496_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_550_inst_ack_0 : boolean;
  signal STORE_col_high_323_store_0_req_1 : boolean;
  signal type_cast_590_inst_req_0 : boolean;
  signal STORE_col_high_323_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_327_inst_req_0 : boolean;
  signal type_cast_623_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_327_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_327_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_327_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_586_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_586_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_550_inst_req_0 : boolean;
  signal STORE_depth_high_329_store_0_req_0 : boolean;
  signal STORE_depth_high_329_store_0_ack_0 : boolean;
  signal STORE_depth_high_329_store_0_req_1 : boolean;
  signal STORE_depth_high_329_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_586_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_586_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_333_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_333_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_333_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_333_inst_ack_1 : boolean;
  signal type_cast_572_inst_ack_1 : boolean;
  signal STORE_pad_335_store_0_req_0 : boolean;
  signal type_cast_572_inst_req_1 : boolean;
  signal STORE_pad_335_store_0_ack_0 : boolean;
  signal STORE_pad_335_store_0_req_1 : boolean;
  signal STORE_pad_335_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_339_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_339_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_514_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_339_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_339_inst_ack_1 : boolean;
  signal type_cast_572_inst_ack_0 : boolean;
  signal type_cast_572_inst_req_0 : boolean;
  signal STORE_out_row_high_341_store_0_req_0 : boolean;
  signal STORE_out_row_high_341_store_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_514_inst_req_1 : boolean;
  signal STORE_out_row_high_341_store_0_req_1 : boolean;
  signal STORE_out_row_high_341_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_345_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_345_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_345_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_345_inst_ack_1 : boolean;
  signal STORE_out_col_high_347_store_0_req_0 : boolean;
  signal STORE_out_col_high_347_store_0_ack_0 : boolean;
  signal type_cast_536_inst_ack_1 : boolean;
  signal STORE_out_col_high_347_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_568_inst_ack_1 : boolean;
  signal STORE_out_col_high_347_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_568_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_351_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_351_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_514_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_351_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_351_inst_ack_1 : boolean;
  signal type_cast_455_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_568_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_568_inst_req_0 : boolean;
  signal type_cast_536_inst_req_1 : boolean;
  signal STORE_out_depth_high_353_store_0_req_0 : boolean;
  signal STORE_out_depth_high_353_store_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_514_inst_req_0 : boolean;
  signal STORE_out_depth_high_353_store_0_req_1 : boolean;
  signal type_cast_554_inst_ack_1 : boolean;
  signal STORE_out_depth_high_353_store_0_ack_1 : boolean;
  signal type_cast_554_inst_req_1 : boolean;
  signal type_cast_554_inst_ack_0 : boolean;
  signal type_cast_554_inst_req_0 : boolean;
  signal LOAD_row_high_357_load_0_req_0 : boolean;
  signal LOAD_row_high_357_load_0_ack_0 : boolean;
  signal LOAD_row_high_357_load_0_req_1 : boolean;
  signal LOAD_row_high_357_load_0_ack_1 : boolean;
  signal type_cast_361_inst_req_0 : boolean;
  signal type_cast_361_inst_ack_0 : boolean;
  signal type_cast_361_inst_req_1 : boolean;
  signal type_cast_361_inst_ack_1 : boolean;
  signal LOAD_col_high_364_load_0_req_0 : boolean;
  signal LOAD_col_high_364_load_0_ack_0 : boolean;
  signal LOAD_col_high_364_load_0_req_1 : boolean;
  signal LOAD_col_high_364_load_0_ack_1 : boolean;
  signal type_cast_368_inst_req_0 : boolean;
  signal type_cast_368_inst_ack_0 : boolean;
  signal type_cast_368_inst_req_1 : boolean;
  signal type_cast_368_inst_ack_1 : boolean;
  signal LOAD_depth_high_371_load_0_req_0 : boolean;
  signal LOAD_depth_high_371_load_0_ack_0 : boolean;
  signal LOAD_depth_high_371_load_0_req_1 : boolean;
  signal LOAD_depth_high_371_load_0_ack_1 : boolean;
  signal type_cast_375_inst_req_0 : boolean;
  signal type_cast_375_inst_ack_0 : boolean;
  signal type_cast_375_inst_req_1 : boolean;
  signal type_cast_375_inst_ack_1 : boolean;
  signal if_stmt_399_branch_req_0 : boolean;
  signal if_stmt_399_branch_ack_1 : boolean;
  signal if_stmt_399_branch_ack_0 : boolean;
  signal type_cast_408_inst_req_0 : boolean;
  signal type_cast_408_inst_ack_0 : boolean;
  signal type_cast_408_inst_req_1 : boolean;
  signal type_cast_408_inst_ack_1 : boolean;
  signal type_cast_412_inst_req_0 : boolean;
  signal type_cast_412_inst_ack_0 : boolean;
  signal type_cast_412_inst_req_1 : boolean;
  signal type_cast_412_inst_ack_1 : boolean;
  signal type_cast_421_inst_req_0 : boolean;
  signal type_cast_421_inst_ack_0 : boolean;
  signal type_cast_421_inst_req_1 : boolean;
  signal type_cast_421_inst_ack_1 : boolean;
  signal array_obj_ref_461_index_offset_req_0 : boolean;
  signal array_obj_ref_461_index_offset_ack_0 : boolean;
  signal array_obj_ref_461_index_offset_req_1 : boolean;
  signal array_obj_ref_461_index_offset_ack_1 : boolean;
  signal addr_of_462_final_reg_req_0 : boolean;
  signal addr_of_462_final_reg_ack_0 : boolean;
  signal addr_of_462_final_reg_req_1 : boolean;
  signal addr_of_462_final_reg_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_465_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_465_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_465_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_465_inst_ack_1 : boolean;
  signal type_cast_469_inst_req_0 : boolean;
  signal type_cast_469_inst_ack_0 : boolean;
  signal type_cast_469_inst_req_1 : boolean;
  signal type_cast_469_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_478_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_478_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_478_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_478_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_689_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_689_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_689_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_689_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_689: Block -- control-path 
    signal testConfigure_CP_689_elements: BooleanArray(132 downto 0);
    -- 
  begin -- 
    testConfigure_CP_689_elements(0) <= testConfigure_CP_689_start;
    testConfigure_CP_689_symbol <= testConfigure_CP_689_elements(125);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	51 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	54 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	66 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	46 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	14 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	19 
    -- CP-element group 0:  members (165) 
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398__entry__
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/ptr_deref_276_Split/split_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/ptr_deref_276_Split/split_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/ptr_deref_276_Split/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/ptr_deref_276_Split/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_base_address_resized
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_268/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/branch_block_stmt_268__entry__
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_update_start_
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_Update/cr
      -- 
    cr_798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => type_cast_285_inst_req_1); -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => STORE_row_high_317_store_0_req_1); -- 
    rr_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => RPIPE_zeropad_input_pipe_281_inst_req_0); -- 
    cr_770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => ptr_deref_276_store_0_req_1); -- 
    cr_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => ptr_deref_294_store_0_req_1); -- 
    cr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => ptr_deref_311_store_0_req_1); -- 
    rr_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => ptr_deref_276_store_0_req_0); -- 
    cr_876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => type_cast_302_inst_req_1); -- 
    cr_1020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => STORE_col_high_323_store_0_req_1); -- 
    cr_1067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => STORE_depth_high_329_store_0_req_1); -- 
    cr_1114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => STORE_pad_335_store_0_req_1); -- 
    cr_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => STORE_out_row_high_341_store_0_req_1); -- 
    cr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => STORE_out_col_high_347_store_0_req_1); -- 
    cr_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => STORE_out_depth_high_353_store_0_req_1); -- 
    cr_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => LOAD_row_high_357_load_0_req_1); -- 
    cr_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => type_cast_361_inst_req_1); -- 
    cr_1330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => LOAD_col_high_364_load_0_req_1); -- 
    cr_1349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => type_cast_368_inst_req_1); -- 
    cr_1377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => LOAD_depth_high_371_load_0_req_1); -- 
    cr_1396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(0), ack => type_cast_375_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	69 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Sample/$exit
      -- 
    ra_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_276_store_0_ack_0, ack => testConfigure_CP_689_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	72 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_Update/$exit
      -- 
    ca_771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_276_store_0_ack_1, ack => testConfigure_CP_689_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_update_start_
      -- CP-element group 3: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_sample_completed_
      -- 
    ra_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_281_inst_ack_0, ack => testConfigure_CP_689_elements(3)); -- 
    cr_784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(3), ack => RPIPE_zeropad_input_pipe_281_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_281_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_Sample/$entry
      -- 
    ca_785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_281_inst_ack_1, ack => testConfigure_CP_689_elements(4)); -- 
    rr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(4), ack => type_cast_285_inst_req_0); -- 
    rr_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(4), ack => RPIPE_zeropad_input_pipe_298_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_Sample/$exit
      -- 
    ra_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_0, ack => testConfigure_CP_689_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_285_update_completed_
      -- 
    ca_799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_1, ack => testConfigure_CP_689_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: 	69 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/word_access_start/$entry
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/word_access_start/word_0/rr
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/ptr_deref_294_Split/split_ack
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/ptr_deref_294_Split/split_req
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/ptr_deref_294_Split/$exit
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/ptr_deref_294_Split/$entry
      -- CP-element group 7: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/$entry
      -- 
    rr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(7), ack => ptr_deref_294_store_0_req_0); -- 
    testConfigure_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(69) & testConfigure_CP_689_elements(6);
      gj_testConfigure_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	70 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/word_access_start/$exit
      -- CP-element group 8: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_sample_completed_
      -- 
    ra_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_294_store_0_ack_0, ack => testConfigure_CP_689_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	72 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_update_completed_
      -- 
    ca_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_294_store_0_ack_1, ack => testConfigure_CP_689_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_update_start_
      -- 
    ra_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_298_inst_ack_0, ack => testConfigure_CP_689_elements(10)); -- 
    cr_862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(10), ack => RPIPE_zeropad_input_pipe_298_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_298_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_Sample/$entry
      -- 
    ca_863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_298_inst_ack_1, ack => testConfigure_CP_689_elements(11)); -- 
    rr_871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(11), ack => type_cast_302_inst_req_0); -- 
    rr_935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(11), ack => RPIPE_zeropad_input_pipe_315_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_Sample/$exit
      -- 
    ra_872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_0, ack => testConfigure_CP_689_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_302_update_completed_
      -- 
    ca_877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_1, ack => testConfigure_CP_689_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	0 
    -- CP-element group 14: 	70 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/ptr_deref_311_Split/split_req
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/ptr_deref_311_Split/$exit
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/ptr_deref_311_Split/$entry
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/word_access_start/word_0/rr
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/ptr_deref_311_Split/split_ack
      -- 
    rr_915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(14), ack => ptr_deref_311_store_0_req_0); -- 
    testConfigure_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(70) & testConfigure_CP_689_elements(13);
      gj_testConfigure_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Sample/word_access_start/$exit
      -- 
    ra_916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_311_store_0_ack_0, ack => testConfigure_CP_689_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	72 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_311_update_completed_
      -- 
    ca_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_311_store_0_ack_1, ack => testConfigure_CP_689_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_update_start_
      -- CP-element group 17: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_sample_completed_
      -- 
    ra_936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_315_inst_ack_0, ack => testConfigure_CP_689_elements(17)); -- 
    cr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(17), ack => RPIPE_zeropad_input_pipe_315_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_315_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_Sample/$entry
      -- 
    ca_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_315_inst_ack_1, ack => testConfigure_CP_689_elements(18)); -- 
    rr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(18), ack => RPIPE_zeropad_input_pipe_321_inst_req_0); -- 
    -- CP-element group 19:  join  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/STORE_row_high_317_Split/$entry
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/word_access_start/word_0/rr
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/word_access_start/$entry
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/STORE_row_high_317_Split/split_ack
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/STORE_row_high_317_Split/split_req
      -- CP-element group 19: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/STORE_row_high_317_Split/$exit
      -- 
    rr_962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(19), ack => STORE_row_high_317_store_0_req_0); -- 
    testConfigure_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(18);
      gj_testConfigure_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	71 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/word_access_start/word_0/ra
      -- CP-element group 20: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Sample/word_access_start/$exit
      -- 
    ra_963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_317_store_0_ack_0, ack => testConfigure_CP_689_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	72 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_Update/$exit
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_317_store_0_ack_1, ack => testConfigure_CP_689_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_update_start_
      -- CP-element group 22: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_Sample/$exit
      -- 
    ra_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_321_inst_ack_0, ack => testConfigure_CP_689_elements(22)); -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(22), ack => RPIPE_zeropad_input_pipe_321_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	27 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_321_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_Sample/rr
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_321_inst_ack_1, ack => testConfigure_CP_689_elements(23)); -- 
    rr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(23), ack => RPIPE_zeropad_input_pipe_327_inst_req_0); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/STORE_col_high_323_Split/$entry
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/STORE_col_high_323_Split/$exit
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/word_access_start/word_0/rr
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/word_access_start/word_0/$entry
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/STORE_col_high_323_Split/split_req
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/STORE_col_high_323_Split/split_ack
      -- CP-element group 24: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/word_access_start/$entry
      -- 
    rr_1009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(24), ack => STORE_col_high_323_store_0_req_0); -- 
    testConfigure_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(23);
      gj_testConfigure_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	67 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_sample_completed_
      -- 
    ra_1010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_323_store_0_ack_0, ack => testConfigure_CP_689_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	72 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_Update/word_access_complete/word_0/ca
      -- 
    ca_1021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_323_store_0_ack_1, ack => testConfigure_CP_689_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_update_start_
      -- CP-element group 27: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_Update/cr
      -- 
    ra_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_327_inst_ack_0, ack => testConfigure_CP_689_elements(27)); -- 
    cr_1034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(27), ack => RPIPE_zeropad_input_pipe_327_inst_req_1); -- 
    -- CP-element group 28:  fork  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	32 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_327_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_Sample/rr
      -- 
    ca_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_327_inst_ack_1, ack => testConfigure_CP_689_elements(28)); -- 
    rr_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(28), ack => RPIPE_zeropad_input_pipe_333_inst_req_0); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (9) 
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/STORE_depth_high_329_Split/$entry
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/STORE_depth_high_329_Split/$exit
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/STORE_depth_high_329_Split/split_req
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/STORE_depth_high_329_Split/split_ack
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/word_access_start/$entry
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/word_access_start/word_0/$entry
      -- CP-element group 29: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/word_access_start/word_0/rr
      -- 
    rr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(29), ack => STORE_depth_high_329_store_0_req_0); -- 
    testConfigure_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(28);
      gj_testConfigure_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	68 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/word_access_start/$exit
      -- CP-element group 30: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/word_access_start/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Sample/word_access_start/word_0/ra
      -- 
    ra_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_329_store_0_ack_0, ack => testConfigure_CP_689_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	72 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Update/word_access_complete/$exit
      -- CP-element group 31: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Update/word_access_complete/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_Update/word_access_complete/word_0/ca
      -- 
    ca_1068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_329_store_0_ack_1, ack => testConfigure_CP_689_elements(31)); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	28 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_update_start_
      -- CP-element group 32: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_Update/cr
      -- 
    ra_1077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_333_inst_ack_0, ack => testConfigure_CP_689_elements(32)); -- 
    cr_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(32), ack => RPIPE_zeropad_input_pipe_333_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: 	37 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_333_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_Sample/rr
      -- 
    ca_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_333_inst_ack_1, ack => testConfigure_CP_689_elements(33)); -- 
    rr_1123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(33), ack => RPIPE_zeropad_input_pipe_339_inst_req_0); -- 
    -- CP-element group 34:  join  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/STORE_pad_335_Split/$entry
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/STORE_pad_335_Split/$exit
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/STORE_pad_335_Split/split_req
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/STORE_pad_335_Split/split_ack
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/word_access_start/$entry
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/word_access_start/word_0/rr
      -- 
    rr_1103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(34), ack => STORE_pad_335_store_0_req_0); -- 
    testConfigure_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(33);
      gj_testConfigure_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/word_access_start/$exit
      -- CP-element group 35: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Sample/word_access_start/word_0/ra
      -- 
    ra_1104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_335_store_0_ack_0, ack => testConfigure_CP_689_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	72 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Update/word_access_complete/$exit
      -- CP-element group 36: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_pad_335_Update/word_access_complete/word_0/ca
      -- 
    ca_1115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_335_store_0_ack_1, ack => testConfigure_CP_689_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	33 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_update_start_
      -- CP-element group 37: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_Update/cr
      -- 
    ra_1124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_339_inst_ack_0, ack => testConfigure_CP_689_elements(37)); -- 
    cr_1128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(37), ack => RPIPE_zeropad_input_pipe_339_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	42 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_339_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_Sample/rr
      -- 
    ca_1129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_339_inst_ack_1, ack => testConfigure_CP_689_elements(38)); -- 
    rr_1170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(38), ack => RPIPE_zeropad_input_pipe_345_inst_req_0); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/STORE_out_row_high_341_Split/$entry
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/STORE_out_row_high_341_Split/$exit
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/STORE_out_row_high_341_Split/split_req
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/STORE_out_row_high_341_Split/split_ack
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/word_access_start/word_0/rr
      -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(39), ack => STORE_out_row_high_341_store_0_req_0); -- 
    testConfigure_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(38);
      gj_testConfigure_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Sample/word_access_start/word_0/ra
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_out_row_high_341_store_0_ack_0, ack => testConfigure_CP_689_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	72 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_row_high_341_Update/word_access_complete/word_0/ca
      -- 
    ca_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_out_row_high_341_store_0_ack_1, ack => testConfigure_CP_689_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	38 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_update_start_
      -- CP-element group 42: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_Update/cr
      -- 
    ra_1171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_345_inst_ack_0, ack => testConfigure_CP_689_elements(42)); -- 
    cr_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(42), ack => RPIPE_zeropad_input_pipe_345_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	47 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_345_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_Sample/rr
      -- 
    ca_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_345_inst_ack_1, ack => testConfigure_CP_689_elements(43)); -- 
    rr_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(43), ack => RPIPE_zeropad_input_pipe_351_inst_req_0); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/STORE_out_col_high_347_Split/$entry
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/STORE_out_col_high_347_Split/$exit
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/STORE_out_col_high_347_Split/split_req
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/STORE_out_col_high_347_Split/split_ack
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/word_access_start/word_0/rr
      -- 
    rr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(44), ack => STORE_out_col_high_347_store_0_req_0); -- 
    testConfigure_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(43);
      gj_testConfigure_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Sample/word_access_start/word_0/ra
      -- 
    ra_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_out_col_high_347_store_0_ack_0, ack => testConfigure_CP_689_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	0 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	72 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_col_high_347_Update/word_access_complete/word_0/ca
      -- 
    ca_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_out_col_high_347_store_0_ack_1, ack => testConfigure_CP_689_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	43 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_update_start_
      -- CP-element group 47: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_Update/cr
      -- 
    ra_1218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_351_inst_ack_0, ack => testConfigure_CP_689_elements(47)); -- 
    cr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(47), ack => RPIPE_zeropad_input_pipe_351_inst_req_1); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/RPIPE_zeropad_input_pipe_351_Update/ca
      -- 
    ca_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_351_inst_ack_1, ack => testConfigure_CP_689_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/STORE_out_depth_high_353_Split/$entry
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/STORE_out_depth_high_353_Split/$exit
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/STORE_out_depth_high_353_Split/split_req
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/STORE_out_depth_high_353_Split/split_ack
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/word_access_start/$entry
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/word_access_start/word_0/$entry
      -- CP-element group 49: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/word_access_start/word_0/rr
      -- 
    rr_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(49), ack => STORE_out_depth_high_353_store_0_req_0); -- 
    testConfigure_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(48);
      gj_testConfigure_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/word_access_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Sample/word_access_start/word_0/ra
      -- 
    ra_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_out_depth_high_353_store_0_ack_0, ack => testConfigure_CP_689_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	0 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	72 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Update/word_access_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_out_depth_high_353_Update/word_access_complete/word_0/ca
      -- 
    ca_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_out_depth_high_353_store_0_ack_1, ack => testConfigure_CP_689_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: 	71 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Sample/word_access_start/$entry
      -- CP-element group 52: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Sample/word_access_start/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Sample/word_access_start/word_0/rr
      -- 
    rr_1272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(52), ack => LOAD_row_high_357_load_0_req_0); -- 
    testConfigure_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(71);
      gj_testConfigure_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Sample/word_access_start/$exit
      -- CP-element group 53: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Sample/word_access_start/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Sample/word_access_start/word_0/ra
      -- 
    ra_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_357_load_0_ack_0, ack => testConfigure_CP_689_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (12) 
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/word_access_complete/$exit
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/word_access_complete/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/word_access_complete/word_0/ca
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/LOAD_row_high_357_Merge/$entry
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/LOAD_row_high_357_Merge/$exit
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/LOAD_row_high_357_Merge/merge_req
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_row_high_357_Update/LOAD_row_high_357_Merge/merge_ack
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_Sample/rr
      -- 
    ca_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_357_load_0_ack_1, ack => testConfigure_CP_689_elements(54)); -- 
    rr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(54), ack => type_cast_361_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_Sample/ra
      -- 
    ra_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_361_inst_ack_0, ack => testConfigure_CP_689_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	72 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_361_Update/ca
      -- 
    ca_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_361_inst_ack_1, ack => testConfigure_CP_689_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: 	67 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Sample/word_access_start/$entry
      -- CP-element group 57: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Sample/word_access_start/word_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Sample/word_access_start/word_0/rr
      -- 
    rr_1319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(57), ack => LOAD_col_high_364_load_0_req_0); -- 
    testConfigure_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(67);
      gj_testConfigure_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (5) 
      -- CP-element group 58: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Sample/word_access_start/$exit
      -- CP-element group 58: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Sample/word_access_start/word_0/$exit
      -- CP-element group 58: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Sample/word_access_start/word_0/ra
      -- 
    ra_1320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_364_load_0_ack_0, ack => testConfigure_CP_689_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (12) 
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/word_access_complete/$exit
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/word_access_complete/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/word_access_complete/word_0/ca
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/LOAD_col_high_364_Merge/$entry
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/LOAD_col_high_364_Merge/$exit
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/LOAD_col_high_364_Merge/merge_req
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_col_high_364_Update/LOAD_col_high_364_Merge/merge_ack
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_Sample/rr
      -- 
    ca_1331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_364_load_0_ack_1, ack => testConfigure_CP_689_elements(59)); -- 
    rr_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(59), ack => type_cast_368_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_Sample/ra
      -- 
    ra_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_368_inst_ack_0, ack => testConfigure_CP_689_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	72 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_368_Update/ca
      -- 
    ca_1350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_368_inst_ack_1, ack => testConfigure_CP_689_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: 	68 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Sample/word_access_start/word_0/rr
      -- 
    rr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(62), ack => LOAD_depth_high_371_load_0_req_0); -- 
    testConfigure_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(0) & testConfigure_CP_689_elements(68);
      gj_testConfigure_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Sample/word_access_start/word_0/ra
      -- 
    ra_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_371_load_0_ack_0, ack => testConfigure_CP_689_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (12) 
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/LOAD_depth_high_371_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/LOAD_depth_high_371_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/LOAD_depth_high_371_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/LOAD_depth_high_371_Update/LOAD_depth_high_371_Merge/merge_ack
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_Sample/rr
      -- 
    ca_1378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_371_load_0_ack_1, ack => testConfigure_CP_689_elements(64)); -- 
    rr_1391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(64), ack => type_cast_375_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_Sample/ra
      -- 
    ra_1392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_375_inst_ack_0, ack => testConfigure_CP_689_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	0 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	72 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/type_cast_375_Update/ca
      -- 
    ca_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_375_inst_ack_1, ack => testConfigure_CP_689_elements(66)); -- 
    -- CP-element group 67:  transition  delay-element  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	57 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_col_high_323_LOAD_col_high_364_delay
      -- 
    -- Element group testConfigure_CP_689_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => testConfigure_CP_689_elements(25), ack => testConfigure_CP_689_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  transition  delay-element  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	30 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	62 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_depth_high_329_LOAD_depth_high_371_delay
      -- 
    -- Element group testConfigure_CP_689_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => testConfigure_CP_689_elements(30), ack => testConfigure_CP_689_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  transition  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	1 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	7 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_276_ptr_deref_294_delay
      -- 
    -- Element group testConfigure_CP_689_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => testConfigure_CP_689_elements(1), ack => testConfigure_CP_689_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  transition  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	8 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	14 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/ptr_deref_294_ptr_deref_311_delay
      -- 
    -- Element group testConfigure_CP_689_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => testConfigure_CP_689_elements(8), ack => testConfigure_CP_689_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  transition  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	20 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	52 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/STORE_row_high_317_LOAD_row_high_357_delay
      -- 
    -- Element group testConfigure_CP_689_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => testConfigure_CP_689_elements(20), ack => testConfigure_CP_689_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  branch  join  transition  place  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	21 
    -- CP-element group 72: 	51 
    -- CP-element group 72: 	56 
    -- CP-element group 72: 	61 
    -- CP-element group 72: 	26 
    -- CP-element group 72: 	66 
    -- CP-element group 72: 	31 
    -- CP-element group 72: 	36 
    -- CP-element group 72: 	41 
    -- CP-element group 72: 	46 
    -- CP-element group 72: 	2 
    -- CP-element group 72: 	9 
    -- CP-element group 72: 	16 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (10) 
      -- CP-element group 72: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398/$exit
      -- CP-element group 72: 	 branch_block_stmt_268/if_stmt_399__entry__
      -- CP-element group 72: 	 branch_block_stmt_268/assign_stmt_274_to_assign_stmt_398__exit__
      -- CP-element group 72: 	 branch_block_stmt_268/if_stmt_399_dead_link/$entry
      -- CP-element group 72: 	 branch_block_stmt_268/if_stmt_399_eval_test/$entry
      -- CP-element group 72: 	 branch_block_stmt_268/if_stmt_399_eval_test/$exit
      -- CP-element group 72: 	 branch_block_stmt_268/if_stmt_399_eval_test/branch_req
      -- CP-element group 72: 	 branch_block_stmt_268/R_cmp72_400_place
      -- CP-element group 72: 	 branch_block_stmt_268/if_stmt_399_if_link/$entry
      -- CP-element group 72: 	 branch_block_stmt_268/if_stmt_399_else_link/$entry
      -- 
    branch_req_1410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(72), ack => if_stmt_399_branch_req_0); -- 
    testConfigure_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(21) & testConfigure_CP_689_elements(51) & testConfigure_CP_689_elements(56) & testConfigure_CP_689_elements(61) & testConfigure_CP_689_elements(26) & testConfigure_CP_689_elements(66) & testConfigure_CP_689_elements(31) & testConfigure_CP_689_elements(36) & testConfigure_CP_689_elements(41) & testConfigure_CP_689_elements(46) & testConfigure_CP_689_elements(2) & testConfigure_CP_689_elements(9) & testConfigure_CP_689_elements(16);
      gj_testConfigure_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  place  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	132 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_268/entry_forx_xend_PhiReq/$exit
      -- CP-element group 73: 	 branch_block_stmt_268/entry_forx_xend_PhiReq/$entry
      -- CP-element group 73: 	 branch_block_stmt_268/if_stmt_399_if_link/$exit
      -- CP-element group 73: 	 branch_block_stmt_268/if_stmt_399_if_link/if_choice_transition
      -- CP-element group 73: 	 branch_block_stmt_268/entry_forx_xend
      -- 
    if_choice_transition_1415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_399_branch_ack_1, ack => testConfigure_CP_689_elements(73)); -- 
    -- CP-element group 74:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74: 	77 
    -- CP-element group 74: 	78 
    -- CP-element group 74: 	79 
    -- CP-element group 74: 	80 
    -- CP-element group 74:  members (30) 
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446__entry__
      -- CP-element group 74: 	 branch_block_stmt_268/merge_stmt_405__exit__
      -- CP-element group 74: 	 branch_block_stmt_268/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_268/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/merge_stmt_405_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_268/merge_stmt_405_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/merge_stmt_405_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_268/merge_stmt_405_PhiAck/dummy
      -- CP-element group 74: 	 branch_block_stmt_268/if_stmt_399_else_link/$exit
      -- CP-element group 74: 	 branch_block_stmt_268/if_stmt_399_else_link/else_choice_transition
      -- CP-element group 74: 	 branch_block_stmt_268/entry_bbx_xnph
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_update_start_
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_update_start_
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_update_start_
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_Update/cr
      -- 
    else_choice_transition_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_399_branch_ack_0, ack => testConfigure_CP_689_elements(74)); -- 
    rr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(74), ack => type_cast_408_inst_req_0); -- 
    cr_1437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(74), ack => type_cast_408_inst_req_1); -- 
    rr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(74), ack => type_cast_412_inst_req_0); -- 
    cr_1451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(74), ack => type_cast_412_inst_req_1); -- 
    rr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(74), ack => type_cast_421_inst_req_0); -- 
    cr_1465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(74), ack => type_cast_421_inst_req_1); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_Sample/ra
      -- 
    ra_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_0, ack => testConfigure_CP_689_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_408_Update/ca
      -- 
    ca_1438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_1, ack => testConfigure_CP_689_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	74 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_Sample/ra
      -- 
    ra_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_412_inst_ack_0, ack => testConfigure_CP_689_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	74 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	81 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_412_Update/ca
      -- 
    ca_1452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_412_inst_ack_1, ack => testConfigure_CP_689_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	74 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_Sample/ra
      -- 
    ra_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_421_inst_ack_0, ack => testConfigure_CP_689_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	74 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/type_cast_421_Update/ca
      -- 
    ca_1466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_421_inst_ack_1, ack => testConfigure_CP_689_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	78 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	126 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_268/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_268/bbx_xnph_forx_xbody
      -- CP-element group 81: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446__exit__
      -- CP-element group 81: 	 branch_block_stmt_268/bbx_xnph_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/$entry
      -- CP-element group 81: 	 branch_block_stmt_268/bbx_xnph_forx_xbody_PhiReq/phi_stmt_449/$entry
      -- CP-element group 81: 	 branch_block_stmt_268/assign_stmt_409_to_assign_stmt_446/$exit
      -- 
    testConfigure_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(76) & testConfigure_CP_689_elements(78) & testConfigure_CP_689_elements(80);
      gj_testConfigure_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	131 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	121 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_sample_complete
      -- CP-element group 82: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_Sample/ack
      -- 
    ack_1495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_461_index_offset_ack_0, ack => testConfigure_CP_689_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	131 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (11) 
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_root_address_calculated
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_offset_calculated
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_Update/ack
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_base_plus_offset/$entry
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_base_plus_offset/$exit
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_base_plus_offset/sum_rename_req
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_base_plus_offset/sum_rename_ack
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_request/$entry
      -- CP-element group 83: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_request/req
      -- 
    ack_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_461_index_offset_ack_1, ack => testConfigure_CP_689_elements(83)); -- 
    req_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(83), ack => addr_of_462_final_reg_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_request/$exit
      -- CP-element group 84: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_request/ack
      -- 
    ack_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_462_final_reg_ack_0, ack => testConfigure_CP_689_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	131 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (19) 
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_addr_resize/$entry
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_addr_resize/$exit
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_addr_resize/base_resize_req
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_root_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_addr_resize/base_resize_ack
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_plus_offset/$entry
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_plus_offset/$exit
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_plus_offset/sum_rename_req
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_plus_offset/sum_rename_ack
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_word_addrgen/$entry
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_word_addrgen/$exit
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_base_address_resized
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_word_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_word_addrgen/root_register_req
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_word_addrgen/root_register_ack
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_complete/$exit
      -- CP-element group 85: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_complete/ack
      -- 
    ack_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_462_final_reg_ack_1, ack => testConfigure_CP_689_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	131 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_update_start_
      -- CP-element group 86: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_Update/cr
      -- 
    ra_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_465_inst_ack_0, ack => testConfigure_CP_689_elements(86)); -- 
    cr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(86), ack => RPIPE_zeropad_input_pipe_465_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_Sample/rr
      -- 
    ca_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_465_inst_ack_1, ack => testConfigure_CP_689_elements(87)); -- 
    rr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(87), ack => type_cast_469_inst_req_0); -- 
    rr_1551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(87), ack => RPIPE_zeropad_input_pipe_478_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_Sample/ra
      -- 
    ra_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_469_inst_ack_0, ack => testConfigure_CP_689_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	131 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_Update/ca
      -- 
    ca_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_469_inst_ack_1, ack => testConfigure_CP_689_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_update_start_
      -- CP-element group 90: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_Update/cr
      -- 
    ra_1552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_478_inst_ack_0, ack => testConfigure_CP_689_elements(90)); -- 
    cr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(90), ack => RPIPE_zeropad_input_pipe_478_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_478_Update/ca
      -- 
    ca_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_478_inst_ack_1, ack => testConfigure_CP_689_elements(91)); -- 
    rr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(91), ack => type_cast_482_inst_req_0); -- 
    rr_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(91), ack => RPIPE_zeropad_input_pipe_496_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_Sample/$exit
      -- 
    ra_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_482_inst_ack_0, ack => testConfigure_CP_689_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	131 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_Update/ca
      -- 
    ca_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_482_inst_ack_1, ack => testConfigure_CP_689_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_update_start_
      -- CP-element group 94: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_Update/cr
      -- 
    ra_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_496_inst_ack_0, ack => testConfigure_CP_689_elements(94)); -- 
    cr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(94), ack => RPIPE_zeropad_input_pipe_496_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_496_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_sample_start_
      -- 
    ca_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_496_inst_ack_1, ack => testConfigure_CP_689_elements(95)); -- 
    rr_1593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(95), ack => type_cast_500_inst_req_0); -- 
    rr_1607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(95), ack => RPIPE_zeropad_input_pipe_514_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_sample_completed_
      -- 
    ra_1594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_500_inst_ack_0, ack => testConfigure_CP_689_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	131 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_Update/ca
      -- 
    ca_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_500_inst_ack_1, ack => testConfigure_CP_689_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_update_start_
      -- CP-element group 98: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_Sample/ra
      -- 
    ra_1608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_514_inst_ack_0, ack => testConfigure_CP_689_elements(98)); -- 
    cr_1612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(98), ack => RPIPE_zeropad_input_pipe_514_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_514_Update/$exit
      -- 
    ca_1613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_514_inst_ack_1, ack => testConfigure_CP_689_elements(99)); -- 
    rr_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(99), ack => type_cast_518_inst_req_0); -- 
    rr_1635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(99), ack => RPIPE_zeropad_input_pipe_532_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_sample_completed_
      -- 
    ra_1622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_0, ack => testConfigure_CP_689_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	131 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_update_completed_
      -- 
    ca_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_1, ack => testConfigure_CP_689_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_update_start_
      -- CP-element group 102: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_Update/cr
      -- 
    ra_1636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_532_inst_ack_0, ack => testConfigure_CP_689_elements(102)); -- 
    cr_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(102), ack => RPIPE_zeropad_input_pipe_532_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_532_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_sample_start_
      -- 
    ca_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_532_inst_ack_1, ack => testConfigure_CP_689_elements(103)); -- 
    rr_1649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(103), ack => type_cast_536_inst_req_0); -- 
    rr_1663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(103), ack => RPIPE_zeropad_input_pipe_550_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_Sample/ra
      -- 
    ra_1650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_536_inst_ack_0, ack => testConfigure_CP_689_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	131 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_Update/$exit
      -- 
    ca_1655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_536_inst_ack_1, ack => testConfigure_CP_689_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_update_start_
      -- CP-element group 106: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_sample_completed_
      -- 
    ra_1664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_550_inst_ack_0, ack => testConfigure_CP_689_elements(106)); -- 
    cr_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(106), ack => RPIPE_zeropad_input_pipe_550_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_550_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_Sample/rr
      -- 
    ca_1669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_550_inst_ack_1, ack => testConfigure_CP_689_elements(107)); -- 
    rr_1677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(107), ack => type_cast_554_inst_req_0); -- 
    rr_1691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(107), ack => RPIPE_zeropad_input_pipe_568_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_Sample/$exit
      -- 
    ra_1678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_554_inst_ack_0, ack => testConfigure_CP_689_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	131 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_Update/ca
      -- CP-element group 109: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_Update/$exit
      -- 
    ca_1683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_554_inst_ack_1, ack => testConfigure_CP_689_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_update_start_
      -- CP-element group 110: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_sample_completed_
      -- 
    ra_1692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_568_inst_ack_0, ack => testConfigure_CP_689_elements(110)); -- 
    cr_1696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(110), ack => RPIPE_zeropad_input_pipe_568_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_568_update_completed_
      -- 
    ca_1697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_568_inst_ack_1, ack => testConfigure_CP_689_elements(111)); -- 
    rr_1705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(111), ack => type_cast_572_inst_req_0); -- 
    rr_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(111), ack => RPIPE_zeropad_input_pipe_586_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_sample_completed_
      -- 
    ra_1706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_572_inst_ack_0, ack => testConfigure_CP_689_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	131 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_update_completed_
      -- 
    ca_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_572_inst_ack_1, ack => testConfigure_CP_689_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_update_start_
      -- CP-element group 114: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_sample_completed_
      -- 
    ra_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_586_inst_ack_0, ack => testConfigure_CP_689_elements(114)); -- 
    cr_1724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(114), ack => RPIPE_zeropad_input_pipe_586_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_586_update_completed_
      -- 
    ca_1725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_586_inst_ack_1, ack => testConfigure_CP_689_elements(115)); -- 
    rr_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(115), ack => type_cast_590_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_sample_completed_
      -- 
    ra_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_590_inst_ack_0, ack => testConfigure_CP_689_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	131 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_update_completed_
      -- 
    ca_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_590_inst_ack_1, ack => testConfigure_CP_689_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/ptr_deref_598_Split/$entry
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/ptr_deref_598_Split/$exit
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/ptr_deref_598_Split/split_req
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/ptr_deref_598_Split/split_ack
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/word_access_start/$entry
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/word_access_start/word_0/$entry
      -- CP-element group 118: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/word_access_start/word_0/rr
      -- 
    rr_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(118), ack => ptr_deref_598_store_0_req_0); -- 
    testConfigure_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(93) & testConfigure_CP_689_elements(97) & testConfigure_CP_689_elements(101) & testConfigure_CP_689_elements(105) & testConfigure_CP_689_elements(109) & testConfigure_CP_689_elements(113) & testConfigure_CP_689_elements(117) & testConfigure_CP_689_elements(85) & testConfigure_CP_689_elements(89);
      gj_testConfigure_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Sample/word_access_start/word_0/ra
      -- 
    ra_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_598_store_0_ack_0, ack => testConfigure_CP_689_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	131 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Update/word_access_complete/word_0/$exit
      -- 
    ca_1789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_598_store_0_ack_1, ack => testConfigure_CP_689_elements(120)); -- 
    -- CP-element group 121:  branch  join  transition  place  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: 	82 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (10) 
      -- CP-element group 121: 	 branch_block_stmt_268/if_stmt_612_eval_test/$entry
      -- CP-element group 121: 	 branch_block_stmt_268/if_stmt_612_dead_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_268/if_stmt_612__entry__
      -- CP-element group 121: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611__exit__
      -- CP-element group 121: 	 branch_block_stmt_268/R_exitcond9_613_place
      -- CP-element group 121: 	 branch_block_stmt_268/if_stmt_612_eval_test/$exit
      -- CP-element group 121: 	 branch_block_stmt_268/if_stmt_612_eval_test/branch_req
      -- CP-element group 121: 	 branch_block_stmt_268/if_stmt_612_if_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_268/if_stmt_612_else_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/$exit
      -- 
    branch_req_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(121), ack => if_stmt_612_branch_req_0); -- 
    testConfigure_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(120) & testConfigure_CP_689_elements(82);
      gj_testConfigure_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  merge  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	132 
    -- CP-element group 122:  members (13) 
      -- CP-element group 122: 	 branch_block_stmt_268/forx_xendx_xloopexit_forx_xend
      -- CP-element group 122: 	 branch_block_stmt_268/merge_stmt_618__exit__
      -- CP-element group 122: 	 branch_block_stmt_268/if_stmt_612_if_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_268/if_stmt_612_if_link/if_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_268/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 122: 	 branch_block_stmt_268/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_268/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_268/merge_stmt_618_PhiAck/dummy
      -- CP-element group 122: 	 branch_block_stmt_268/merge_stmt_618_PhiAck/$exit
      -- CP-element group 122: 	 branch_block_stmt_268/merge_stmt_618_PhiAck/$entry
      -- CP-element group 122: 	 branch_block_stmt_268/merge_stmt_618_PhiReqMerge
      -- CP-element group 122: 	 branch_block_stmt_268/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_268/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_612_branch_ack_1, ack => testConfigure_CP_689_elements(122)); -- 
    -- CP-element group 123:  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	127 
    -- CP-element group 123: 	128 
    -- CP-element group 123:  members (12) 
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/$entry
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/Update/cr
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/$entry
      -- CP-element group 123: 	 branch_block_stmt_268/if_stmt_612_else_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/$entry
      -- CP-element group 123: 	 branch_block_stmt_268/if_stmt_612_else_link/else_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/$entry
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_268/forx_xbody_forx_xbody
      -- 
    else_choice_transition_1806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_612_branch_ack_0, ack => testConfigure_CP_689_elements(123)); -- 
    cr_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(123), ack => type_cast_455_inst_req_1); -- 
    rr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(123), ack => type_cast_455_inst_req_0); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	132 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_Sample/ra
      -- CP-element group 124: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_sample_completed_
      -- 
    ra_1820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_0, ack => testConfigure_CP_689_elements(124)); -- 
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	132 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (16) 
      -- CP-element group 125: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_268/merge_stmt_626__exit__
      -- CP-element group 125: 	 branch_block_stmt_268/return__
      -- CP-element group 125: 	 branch_block_stmt_268/branch_block_stmt_268__exit__
      -- CP-element group 125: 	 branch_block_stmt_268/assign_stmt_624__exit__
      -- CP-element group 125: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_268/return___PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_268/return___PhiReq/$exit
      -- CP-element group 125: 	 branch_block_stmt_268/merge_stmt_626_PhiReqMerge
      -- CP-element group 125: 	 branch_block_stmt_268/merge_stmt_626_PhiAck/$entry
      -- CP-element group 125: 	 branch_block_stmt_268/merge_stmt_626_PhiAck/$exit
      -- CP-element group 125: 	 branch_block_stmt_268/merge_stmt_626_PhiAck/dummy
      -- CP-element group 125: 	 $exit
      -- CP-element group 125: 	 branch_block_stmt_268/$exit
      -- CP-element group 125: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_268/assign_stmt_624/$exit
      -- 
    ca_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_1, ack => testConfigure_CP_689_elements(125)); -- 
    -- CP-element group 126:  transition  output  delay-element  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	81 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	130 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_268/bbx_xnph_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_req
      -- CP-element group 126: 	 branch_block_stmt_268/bbx_xnph_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_453_konst_delay_trans
      -- CP-element group 126: 	 branch_block_stmt_268/bbx_xnph_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_268/bbx_xnph_forx_xbody_PhiReq/phi_stmt_449/$exit
      -- CP-element group 126: 	 branch_block_stmt_268/bbx_xnph_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_449_req_1848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_449_req_1848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(126), ack => phi_stmt_449_req_0); -- 
    -- Element group testConfigure_CP_689_elements(126) is a control-delay.
    cp_element_126_delay: control_delay_element  generic map(name => " 126_delay", delay_value => 1)  port map(req => testConfigure_CP_689_elements(81), ack => testConfigure_CP_689_elements(126), clk => clk, reset =>reset);
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	123 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/Sample/ra
      -- 
    ra_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_455_inst_ack_0, ack => testConfigure_CP_689_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	123 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/Update/ca
      -- 
    ca_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_455_inst_ack_1, ack => testConfigure_CP_689_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_req
      -- CP-element group 129: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/$exit
      -- CP-element group 129: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 129: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/phi_stmt_449_sources/type_cast_455/$exit
      -- CP-element group 129: 	 branch_block_stmt_268/forx_xbody_forx_xbody_PhiReq/phi_stmt_449/$exit
      -- 
    phi_stmt_449_req_1874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_449_req_1874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(129), ack => phi_stmt_449_req_1); -- 
    testConfigure_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_689_elements(127) & testConfigure_CP_689_elements(128);
      gj_testConfigure_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_689_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	126 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_268/merge_stmt_448_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_268/merge_stmt_448_PhiAck/$entry
      -- 
    testConfigure_CP_689_elements(130) <= OrReduce(testConfigure_CP_689_elements(126) & testConfigure_CP_689_elements(129));
    -- CP-element group 131:  fork  transition  place  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	93 
    -- CP-element group 131: 	97 
    -- CP-element group 131: 	101 
    -- CP-element group 131: 	105 
    -- CP-element group 131: 	109 
    -- CP-element group 131: 	113 
    -- CP-element group 131: 	117 
    -- CP-element group 131: 	120 
    -- CP-element group 131: 	82 
    -- CP-element group 131: 	83 
    -- CP-element group 131: 	85 
    -- CP-element group 131: 	86 
    -- CP-element group 131: 	89 
    -- CP-element group 131:  members (56) 
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_482_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611__entry__
      -- CP-element group 131: 	 branch_block_stmt_268/merge_stmt_448__exit__
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_500_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/merge_stmt_448_PhiAck/$exit
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Update/word_access_complete/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/merge_stmt_448_PhiAck/phi_stmt_449_ack
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Update/word_access_complete/word_0/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/ptr_deref_598_Update/word_access_complete/word_0/cr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_590_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_518_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_572_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_554_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_536_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_resized_1
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_scaled_1
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_computed_1
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_resize_1/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_resize_1/$exit
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_resize_1/index_resize_req
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_resize_1/index_resize_ack
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_scale_1/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_scale_1/$exit
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_scale_1/scale_rename_req
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_index_scale_1/scale_rename_ack
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_update_start
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_Sample/req
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/array_obj_ref_461_final_index_sum_regn_Update/req
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_complete/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/addr_of_462_complete/req
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/RPIPE_zeropad_input_pipe_465_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_update_start_
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_268/assign_stmt_463_to_assign_stmt_611/type_cast_469_Update/cr
      -- 
    phi_stmt_449_ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_449_ack_0, ack => testConfigure_CP_689_elements(131)); -- 
    cr_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => type_cast_590_inst_req_1); -- 
    cr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => type_cast_482_inst_req_1); -- 
    cr_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => type_cast_518_inst_req_1); -- 
    cr_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => type_cast_500_inst_req_1); -- 
    cr_1788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => ptr_deref_598_store_0_req_1); -- 
    cr_1710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => type_cast_572_inst_req_1); -- 
    cr_1654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => type_cast_536_inst_req_1); -- 
    cr_1682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => type_cast_554_inst_req_1); -- 
    req_1494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => array_obj_ref_461_index_offset_req_0); -- 
    req_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => array_obj_ref_461_index_offset_req_1); -- 
    req_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => addr_of_462_final_reg_req_1); -- 
    rr_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => RPIPE_zeropad_input_pipe_465_inst_req_0); -- 
    cr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(131), ack => type_cast_469_inst_req_1); -- 
    -- CP-element group 132:  merge  fork  transition  place  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	122 
    -- CP-element group 132: 	73 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	124 
    -- CP-element group 132: 	125 
    -- CP-element group 132:  members (13) 
      -- CP-element group 132: 	 branch_block_stmt_268/merge_stmt_620_PhiAck/$entry
      -- CP-element group 132: 	 branch_block_stmt_268/merge_stmt_620_PhiAck/$exit
      -- CP-element group 132: 	 branch_block_stmt_268/merge_stmt_620_PhiAck/dummy
      -- CP-element group 132: 	 branch_block_stmt_268/assign_stmt_624__entry__
      -- CP-element group 132: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_268/merge_stmt_620__exit__
      -- CP-element group 132: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_268/merge_stmt_620_PhiReqMerge
      -- CP-element group 132: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_update_start_
      -- CP-element group 132: 	 branch_block_stmt_268/assign_stmt_624/type_cast_623_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_268/assign_stmt_624/$entry
      -- 
    cr_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(132), ack => type_cast_623_inst_req_1); -- 
    rr_1819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_689_elements(132), ack => type_cast_623_inst_req_0); -- 
    testConfigure_CP_689_elements(132) <= OrReduce(testConfigure_CP_689_elements(122) & testConfigure_CP_689_elements(73));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_col_high_364_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_364_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_371_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_371_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_357_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_357_word_address_0 : std_logic_vector(0 downto 0);
    signal R_indvar_460_resized : std_logic_vector(13 downto 0);
    signal R_indvar_460_scaled : std_logic_vector(13 downto 0);
    signal STORE_col_high_323_data_0 : std_logic_vector(7 downto 0);
    signal STORE_col_high_323_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_depth_high_329_data_0 : std_logic_vector(7 downto 0);
    signal STORE_depth_high_329_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_out_col_high_347_data_0 : std_logic_vector(7 downto 0);
    signal STORE_out_col_high_347_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_out_depth_high_353_data_0 : std_logic_vector(7 downto 0);
    signal STORE_out_depth_high_353_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_out_row_high_341_data_0 : std_logic_vector(7 downto 0);
    signal STORE_out_row_high_341_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_pad_335_data_0 : std_logic_vector(7 downto 0);
    signal STORE_pad_335_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_row_high_317_data_0 : std_logic_vector(7 downto 0);
    signal STORE_row_high_317_word_address_0 : std_logic_vector(0 downto 0);
    signal add33_506 : std_logic_vector(63 downto 0);
    signal add39_524 : std_logic_vector(63 downto 0);
    signal add45_542 : std_logic_vector(63 downto 0);
    signal add51_560 : std_logic_vector(63 downto 0);
    signal add57_578 : std_logic_vector(63 downto 0);
    signal add63_596 : std_logic_vector(63 downto 0);
    signal add_488 : std_logic_vector(63 downto 0);
    signal array_obj_ref_461_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_461_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_461_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_461_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_461_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_461_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_463 : std_logic_vector(31 downto 0);
    signal call1_299 : std_logic_vector(7 downto 0);
    signal call22_466 : std_logic_vector(7 downto 0);
    signal call25_479 : std_logic_vector(7 downto 0);
    signal call30_497 : std_logic_vector(7 downto 0);
    signal call36_515 : std_logic_vector(7 downto 0);
    signal call3_316 : std_logic_vector(7 downto 0);
    signal call42_533 : std_logic_vector(7 downto 0);
    signal call48_551 : std_logic_vector(7 downto 0);
    signal call4_322 : std_logic_vector(7 downto 0);
    signal call54_569 : std_logic_vector(7 downto 0);
    signal call5_328 : std_logic_vector(7 downto 0);
    signal call60_587 : std_logic_vector(7 downto 0);
    signal call6_334 : std_logic_vector(7 downto 0);
    signal call7_340 : std_logic_vector(7 downto 0);
    signal call8_346 : std_logic_vector(7 downto 0);
    signal call9_352 : std_logic_vector(7 downto 0);
    signal call_282 : std_logic_vector(7 downto 0);
    signal cmp72_398 : std_logic_vector(0 downto 0);
    signal conv10_362 : std_logic_vector(63 downto 0);
    signal conv12_369 : std_logic_vector(63 downto 0);
    signal conv14_376 : std_logic_vector(63 downto 0);
    signal conv23_470 : std_logic_vector(63 downto 0);
    signal conv27_483 : std_logic_vector(63 downto 0);
    signal conv2_303 : std_logic_vector(31 downto 0);
    signal conv32_501 : std_logic_vector(63 downto 0);
    signal conv38_519 : std_logic_vector(63 downto 0);
    signal conv44_537 : std_logic_vector(63 downto 0);
    signal conv50_555 : std_logic_vector(63 downto 0);
    signal conv56_573 : std_logic_vector(63 downto 0);
    signal conv62_591 : std_logic_vector(63 downto 0);
    signal conv_286 : std_logic_vector(31 downto 0);
    signal exitcond9_611 : std_logic_vector(0 downto 0);
    signal iNsTr_0_274 : std_logic_vector(31 downto 0);
    signal iNsTr_3_292 : std_logic_vector(31 downto 0);
    signal iNsTr_6_309 : std_logic_vector(31 downto 0);
    signal indvar_449 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_606 : std_logic_vector(63 downto 0);
    signal mul15_386 : std_logic_vector(63 downto 0);
    signal mul_381 : std_logic_vector(63 downto 0);
    signal ptr_deref_276_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_276_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_276_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_276_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_276_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_276_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_294_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_294_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_294_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_294_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_294_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_294_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_311_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_311_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_311_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_311_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_311_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_311_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_598_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_598_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_598_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_598_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_598_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_598_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl29_494 : std_logic_vector(63 downto 0);
    signal shl35_512 : std_logic_vector(63 downto 0);
    signal shl41_530 : std_logic_vector(63 downto 0);
    signal shl47_548 : std_logic_vector(63 downto 0);
    signal shl53_566 : std_logic_vector(63 downto 0);
    signal shl59_584 : std_logic_vector(63 downto 0);
    signal shl_476 : std_logic_vector(63 downto 0);
    signal shr71x_xmask_392 : std_logic_vector(63 downto 0);
    signal tmp11_365 : std_logic_vector(7 downto 0);
    signal tmp13_372 : std_logic_vector(7 downto 0);
    signal tmp1_409 : std_logic_vector(63 downto 0);
    signal tmp2_413 : std_logic_vector(63 downto 0);
    signal tmp3_418 : std_logic_vector(63 downto 0);
    signal tmp4_422 : std_logic_vector(63 downto 0);
    signal tmp5_427 : std_logic_vector(63 downto 0);
    signal tmp6_433 : std_logic_vector(63 downto 0);
    signal tmp7_439 : std_logic_vector(0 downto 0);
    signal tmp_358 : std_logic_vector(7 downto 0);
    signal type_cast_278_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_390_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_396_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_431_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_437_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_444_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_453_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_455_wire : std_logic_vector(63 downto 0);
    signal type_cast_474_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_492_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_510_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_528_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_546_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_564_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_604_wire_constant : std_logic_vector(63 downto 0);
    signal umax8_446 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    LOAD_col_high_364_word_address_0 <= "0";
    LOAD_depth_high_371_word_address_0 <= "0";
    LOAD_row_high_357_word_address_0 <= "0";
    STORE_col_high_323_word_address_0 <= "0";
    STORE_depth_high_329_word_address_0 <= "0";
    STORE_out_col_high_347_word_address_0 <= "0";
    STORE_out_depth_high_353_word_address_0 <= "0";
    STORE_out_row_high_341_word_address_0 <= "0";
    STORE_pad_335_word_address_0 <= "0";
    STORE_row_high_317_word_address_0 <= "0";
    array_obj_ref_461_constant_part_of_offset <= "00000000000000";
    array_obj_ref_461_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_461_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_461_resized_base_address <= "00000000000000";
    iNsTr_0_274 <= "00000000000000000000000000000000";
    iNsTr_3_292 <= "00000000000000000000000000000001";
    iNsTr_6_309 <= "00000000000000000000000000000010";
    ptr_deref_276_word_offset_0 <= "0000000";
    ptr_deref_294_word_offset_0 <= "0000000";
    ptr_deref_311_word_offset_0 <= "0000000";
    ptr_deref_598_word_offset_0 <= "00000000000000";
    type_cast_278_wire_constant <= "00000000000000000000000000000101";
    type_cast_390_wire_constant <= "0000000000000000000000000000000000000000111111111111111111111100";
    type_cast_396_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_431_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_437_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_444_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_453_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_474_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_492_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_510_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_528_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_546_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_564_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_582_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_604_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_449: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_453_wire_constant & type_cast_455_wire;
      req <= phi_stmt_449_req_0 & phi_stmt_449_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_449",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_449_ack_0,
          idata => idata,
          odata => indvar_449,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_449
    -- flow-through select operator MUX_445_inst
    umax8_446 <= tmp6_433 when (tmp7_439(0) /=  '0') else type_cast_444_wire_constant;
    addr_of_462_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_462_final_reg_req_0;
      addr_of_462_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_462_final_reg_req_1;
      addr_of_462_final_reg_ack_1<= rack(0);
      addr_of_462_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_462_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_461_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_463,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_285_inst_req_0;
      type_cast_285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_285_inst_req_1;
      type_cast_285_inst_ack_1<= rack(0);
      type_cast_285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_302_inst_req_0;
      type_cast_302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_302_inst_req_1;
      type_cast_302_inst_ack_1<= rack(0);
      type_cast_302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_361_inst_req_0;
      type_cast_361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_361_inst_req_1;
      type_cast_361_inst_ack_1<= rack(0);
      type_cast_361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_368_inst_req_0;
      type_cast_368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_368_inst_req_1;
      type_cast_368_inst_ack_1<= rack(0);
      type_cast_368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_375_inst_req_0;
      type_cast_375_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_375_inst_req_1;
      type_cast_375_inst_ack_1<= rack(0);
      type_cast_375_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_375_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp13_372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_376,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_408_inst_req_0;
      type_cast_408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_408_inst_req_1;
      type_cast_408_inst_ack_1<= rack(0);
      type_cast_408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_412_inst_req_0;
      type_cast_412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_412_inst_req_1;
      type_cast_412_inst_ack_1<= rack(0);
      type_cast_412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp2_413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_421_inst_req_0;
      type_cast_421_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_421_inst_req_1;
      type_cast_421_inst_ack_1<= rack(0);
      type_cast_421_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_421_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp13_372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp4_422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_455_inst_req_0;
      type_cast_455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_455_inst_req_1;
      type_cast_455_inst_ack_1<= rack(0);
      type_cast_455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_606,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_455_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_469_inst_req_0;
      type_cast_469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_469_inst_req_1;
      type_cast_469_inst_ack_1<= rack(0);
      type_cast_469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_482_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_482_inst_req_0;
      type_cast_482_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_482_inst_req_1;
      type_cast_482_inst_ack_1<= rack(0);
      type_cast_482_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_482_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call25_479,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_500_inst_req_0;
      type_cast_500_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_500_inst_req_1;
      type_cast_500_inst_ack_1<= rack(0);
      type_cast_500_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_500_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call30_497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_501,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_518_inst_req_0;
      type_cast_518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_518_inst_req_1;
      type_cast_518_inst_ack_1<= rack(0);
      type_cast_518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_536_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_536_inst_req_0;
      type_cast_536_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_536_inst_req_1;
      type_cast_536_inst_ack_1<= rack(0);
      type_cast_536_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_536_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_533,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_537,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_554_inst_req_0;
      type_cast_554_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_554_inst_req_1;
      type_cast_554_inst_ack_1<= rack(0);
      type_cast_554_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call48_551,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_555,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_572_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_572_inst_req_0;
      type_cast_572_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_572_inst_req_1;
      type_cast_572_inst_ack_1<= rack(0);
      type_cast_572_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_572_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call54_569,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_573,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_590_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_590_inst_req_0;
      type_cast_590_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_590_inst_req_1;
      type_cast_590_inst_ack_1<= rack(0);
      type_cast_590_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_590_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call60_587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_623_inst_req_0;
      type_cast_623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_623_inst_req_1;
      type_cast_623_inst_ack_1<= rack(0);
      type_cast_623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_623_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul15_386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_col_high_364_gather_scatter
    process(LOAD_col_high_364_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_364_data_0;
      ov(7 downto 0) := iv;
      tmp11_365 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_371_gather_scatter
    process(LOAD_depth_high_371_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_371_data_0;
      ov(7 downto 0) := iv;
      tmp13_372 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_357_gather_scatter
    process(LOAD_row_high_357_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_357_data_0;
      ov(7 downto 0) := iv;
      tmp_358 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_col_high_323_gather_scatter
    process(call4_322) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call4_322;
      ov(7 downto 0) := iv;
      STORE_col_high_323_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_depth_high_329_gather_scatter
    process(call5_328) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call5_328;
      ov(7 downto 0) := iv;
      STORE_depth_high_329_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_out_col_high_347_gather_scatter
    process(call8_346) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call8_346;
      ov(7 downto 0) := iv;
      STORE_out_col_high_347_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_out_depth_high_353_gather_scatter
    process(call9_352) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call9_352;
      ov(7 downto 0) := iv;
      STORE_out_depth_high_353_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_out_row_high_341_gather_scatter
    process(call7_340) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call7_340;
      ov(7 downto 0) := iv;
      STORE_out_row_high_341_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_pad_335_gather_scatter
    process(call6_334) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call6_334;
      ov(7 downto 0) := iv;
      STORE_pad_335_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_row_high_317_gather_scatter
    process(call3_316) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call3_316;
      ov(7 downto 0) := iv;
      STORE_row_high_317_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_461_index_1_rename
    process(R_indvar_460_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_460_resized;
      ov(13 downto 0) := iv;
      R_indvar_460_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_461_index_1_resize
    process(indvar_449) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_449;
      ov := iv(13 downto 0);
      R_indvar_460_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_461_root_address_inst
    process(array_obj_ref_461_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_461_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_461_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_276_addr_0
    process(ptr_deref_276_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_276_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_276_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_276_base_resize
    process(iNsTr_0_274) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_274;
      ov := iv(6 downto 0);
      ptr_deref_276_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_276_gather_scatter
    process(type_cast_278_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_278_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_276_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_276_root_address_inst
    process(ptr_deref_276_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_276_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_276_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_294_addr_0
    process(ptr_deref_294_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_294_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_294_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_294_base_resize
    process(iNsTr_3_292) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_292;
      ov := iv(6 downto 0);
      ptr_deref_294_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_294_gather_scatter
    process(conv_286) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_286;
      ov(31 downto 0) := iv;
      ptr_deref_294_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_294_root_address_inst
    process(ptr_deref_294_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_294_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_294_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_311_addr_0
    process(ptr_deref_311_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_311_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_311_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_311_base_resize
    process(iNsTr_6_309) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_309;
      ov := iv(6 downto 0);
      ptr_deref_311_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_311_gather_scatter
    process(conv2_303) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv2_303;
      ov(31 downto 0) := iv;
      ptr_deref_311_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_311_root_address_inst
    process(ptr_deref_311_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_311_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_311_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_598_addr_0
    process(ptr_deref_598_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_598_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_598_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_598_base_resize
    process(arrayidx_463) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_463;
      ov := iv(13 downto 0);
      ptr_deref_598_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_598_gather_scatter
    process(add63_596) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add63_596;
      ov(63 downto 0) := iv;
      ptr_deref_598_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_598_root_address_inst
    process(ptr_deref_598_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_598_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_598_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_399_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp72_398;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_399_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_399_branch_req_0,
          ack0 => if_stmt_399_branch_ack_0,
          ack1 => if_stmt_399_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_612_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond9_611;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_612_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_612_branch_req_0,
          ack0 => if_stmt_612_branch_ack_0,
          ack1 => if_stmt_612_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_605_inst
    process(indvar_449) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_449, type_cast_604_wire_constant, tmp_var);
      indvarx_xnext_606 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_391_inst
    process(mul15_386) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul15_386, type_cast_390_wire_constant, tmp_var);
      shr71x_xmask_392 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_397_inst
    process(shr71x_xmask_392) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr71x_xmask_392, type_cast_396_wire_constant, tmp_var);
      cmp72_398 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_610_inst
    process(indvarx_xnext_606, umax8_446) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_606, umax8_446, tmp_var);
      exitcond9_611 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_432_inst
    process(tmp5_427) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_427, type_cast_431_wire_constant, tmp_var);
      tmp6_433 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_380_inst
    process(conv12_369, conv10_362) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv12_369, conv10_362, tmp_var);
      mul_381 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_385_inst
    process(mul_381, conv14_376) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_381, conv14_376, tmp_var);
      mul15_386 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_417_inst
    process(tmp1_409, tmp2_413) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_409, tmp2_413, tmp_var);
      tmp3_418 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_426_inst
    process(tmp3_418, tmp4_422) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_418, tmp4_422, tmp_var);
      tmp5_427 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_487_inst
    process(shl_476, conv27_483) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_476, conv27_483, tmp_var);
      add_488 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_505_inst
    process(shl29_494, conv32_501) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl29_494, conv32_501, tmp_var);
      add33_506 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_523_inst
    process(shl35_512, conv38_519) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl35_512, conv38_519, tmp_var);
      add39_524 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_541_inst
    process(shl41_530, conv44_537) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl41_530, conv44_537, tmp_var);
      add45_542 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_559_inst
    process(shl47_548, conv50_555) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl47_548, conv50_555, tmp_var);
      add51_560 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_577_inst
    process(shl53_566, conv56_573) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl53_566, conv56_573, tmp_var);
      add57_578 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_595_inst
    process(shl59_584, conv62_591) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl59_584, conv62_591, tmp_var);
      add63_596 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_475_inst
    process(conv23_470) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv23_470, type_cast_474_wire_constant, tmp_var);
      shl_476 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_493_inst
    process(add_488) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_488, type_cast_492_wire_constant, tmp_var);
      shl29_494 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_511_inst
    process(add33_506) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add33_506, type_cast_510_wire_constant, tmp_var);
      shl35_512 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_529_inst
    process(add39_524) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add39_524, type_cast_528_wire_constant, tmp_var);
      shl41_530 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_547_inst
    process(add45_542) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add45_542, type_cast_546_wire_constant, tmp_var);
      shl47_548 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_565_inst
    process(add51_560) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add51_560, type_cast_564_wire_constant, tmp_var);
      shl53_566 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_583_inst
    process(add57_578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add57_578, type_cast_582_wire_constant, tmp_var);
      shl59_584 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_438_inst
    process(tmp6_433) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp6_433, type_cast_437_wire_constant, tmp_var);
      tmp7_439 <= tmp_var; --
    end process;
    -- shared split operator group (24) : array_obj_ref_461_index_offset 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_460_scaled;
      array_obj_ref_461_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_461_index_offset_req_0;
      array_obj_ref_461_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_461_index_offset_req_1;
      array_obj_ref_461_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared load operator group (0) : LOAD_col_high_364_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_col_high_364_load_0_req_0;
      LOAD_col_high_364_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_col_high_364_load_0_req_1;
      LOAD_col_high_364_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_col_high_364_word_address_0;
      LOAD_col_high_364_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : LOAD_depth_high_371_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_depth_high_371_load_0_req_0;
      LOAD_depth_high_371_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_depth_high_371_load_0_req_1;
      LOAD_depth_high_371_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_depth_high_371_word_address_0;
      LOAD_depth_high_371_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(7 downto 0),
          mtag => memory_space_4_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : LOAD_row_high_357_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_row_high_357_load_0_req_0;
      LOAD_row_high_357_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_row_high_357_load_0_req_1;
      LOAD_row_high_357_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_row_high_357_word_address_0;
      LOAD_row_high_357_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(0),
          mack => memory_space_10_lr_ack(0),
          maddr => memory_space_10_lr_addr(0 downto 0),
          mtag => memory_space_10_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(0),
          mack => memory_space_10_lc_ack(0),
          mdata => memory_space_10_lc_data(7 downto 0),
          mtag => memory_space_10_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : STORE_col_high_323_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_col_high_323_store_0_req_0;
      STORE_col_high_323_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_col_high_323_store_0_req_1;
      STORE_col_high_323_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_col_high_323_word_address_0;
      data_in <= STORE_col_high_323_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : STORE_depth_high_329_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_depth_high_329_store_0_req_0;
      STORE_depth_high_329_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_depth_high_329_store_0_req_1;
      STORE_depth_high_329_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_depth_high_329_word_address_0;
      data_in <= STORE_depth_high_329_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : STORE_out_col_high_347_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_out_col_high_347_store_0_req_0;
      STORE_out_col_high_347_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_out_col_high_347_store_0_req_1;
      STORE_out_col_high_347_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_out_col_high_347_word_address_0;
      data_in <= STORE_out_col_high_347_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(7 downto 0),
          mtag => memory_space_6_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : STORE_out_depth_high_353_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_out_depth_high_353_store_0_req_0;
      STORE_out_depth_high_353_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_out_depth_high_353_store_0_req_1;
      STORE_out_depth_high_353_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_out_depth_high_353_word_address_0;
      data_in <= STORE_out_depth_high_353_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(7 downto 0),
          mtag => memory_space_7_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : STORE_out_row_high_341_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_out_row_high_341_store_0_req_0;
      STORE_out_row_high_341_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_out_row_high_341_store_0_req_1;
      STORE_out_row_high_341_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_out_row_high_341_word_address_0;
      data_in <= STORE_out_row_high_341_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : STORE_pad_335_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_pad_335_store_0_req_0;
      STORE_pad_335_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_pad_335_store_0_req_1;
      STORE_pad_335_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_pad_335_word_address_0;
      data_in <= STORE_pad_335_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_9_sr_req(0),
          mack => memory_space_9_sr_ack(0),
          maddr => memory_space_9_sr_addr(0 downto 0),
          mdata => memory_space_9_sr_data(7 downto 0),
          mtag => memory_space_9_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_9_sc_req(0),
          mack => memory_space_9_sc_ack(0),
          mtag => memory_space_9_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : STORE_row_high_317_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_row_high_317_store_0_req_0;
      STORE_row_high_317_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_row_high_317_store_0_req_1;
      STORE_row_high_317_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_row_high_317_word_address_0;
      data_in <= STORE_row_high_317_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_10_sr_req(0),
          mack => memory_space_10_sr_ack(0),
          maddr => memory_space_10_sr_addr(0 downto 0),
          mdata => memory_space_10_sr_data(7 downto 0),
          mtag => memory_space_10_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_10_sc_req(0),
          mack => memory_space_10_sc_ack(0),
          mtag => memory_space_10_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_276_store_0 ptr_deref_294_store_0 ptr_deref_311_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_276_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_294_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_311_store_0_req_0;
      ptr_deref_276_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_294_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_311_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_276_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_294_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_311_store_0_req_1;
      ptr_deref_276_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_294_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_311_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup7_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup7_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup7_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup7_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup7_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup7_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup7_gI: SplitGuardInterface generic map(name => "StoreGroup7_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_276_word_address_0 & ptr_deref_294_word_address_0 & ptr_deref_311_word_address_0;
      data_in <= ptr_deref_276_data_0 & ptr_deref_294_data_0 & ptr_deref_311_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup7 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(6 downto 0),
          mdata => memory_space_5_sr_data(31 downto 0),
          mtag => memory_space_5_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup7 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared store operator group (8) : ptr_deref_598_store_0 
    StoreGroup8: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_598_store_0_req_0;
      ptr_deref_598_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_598_store_0_req_1;
      ptr_deref_598_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup8_gI: SplitGuardInterface generic map(name => "StoreGroup8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_598_word_address_0;
      data_in <= ptr_deref_598_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup8 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup8 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 8
    -- shared inport operator group (0) : RPIPE_zeropad_input_pipe_281_inst RPIPE_zeropad_input_pipe_298_inst RPIPE_zeropad_input_pipe_315_inst RPIPE_zeropad_input_pipe_321_inst RPIPE_zeropad_input_pipe_327_inst RPIPE_zeropad_input_pipe_333_inst RPIPE_zeropad_input_pipe_339_inst RPIPE_zeropad_input_pipe_345_inst RPIPE_zeropad_input_pipe_351_inst RPIPE_zeropad_input_pipe_465_inst RPIPE_zeropad_input_pipe_478_inst RPIPE_zeropad_input_pipe_496_inst RPIPE_zeropad_input_pipe_514_inst RPIPE_zeropad_input_pipe_532_inst RPIPE_zeropad_input_pipe_550_inst RPIPE_zeropad_input_pipe_568_inst RPIPE_zeropad_input_pipe_586_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(135 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 16 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 16 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 16 downto 0);
      signal guard_vector : std_logic_vector( 16 downto 0);
      constant outBUFs : IntegerArray(16 downto 0) := (16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(16 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false);
      constant guardBuffering: IntegerArray(16 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2);
      -- 
    begin -- 
      reqL_unguarded(16) <= RPIPE_zeropad_input_pipe_281_inst_req_0;
      reqL_unguarded(15) <= RPIPE_zeropad_input_pipe_298_inst_req_0;
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_315_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_321_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_327_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_333_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_339_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_345_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_351_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_465_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_478_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_496_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_514_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_532_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_550_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_568_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_586_inst_req_0;
      RPIPE_zeropad_input_pipe_281_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_zeropad_input_pipe_298_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_zeropad_input_pipe_315_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_321_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_327_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_333_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_339_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_345_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_351_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_465_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_478_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_496_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_514_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_532_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_550_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_568_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_586_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(16) <= RPIPE_zeropad_input_pipe_281_inst_req_1;
      reqR_unguarded(15) <= RPIPE_zeropad_input_pipe_298_inst_req_1;
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_315_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_321_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_327_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_333_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_339_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_345_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_351_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_465_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_478_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_496_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_514_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_532_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_550_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_568_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_586_inst_req_1;
      RPIPE_zeropad_input_pipe_281_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_zeropad_input_pipe_298_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_zeropad_input_pipe_315_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_321_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_327_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_333_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_339_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_345_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_351_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_465_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_478_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_496_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_514_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_532_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_550_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_568_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_586_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      call_282 <= data_out(135 downto 128);
      call1_299 <= data_out(127 downto 120);
      call3_316 <= data_out(119 downto 112);
      call4_322 <= data_out(111 downto 104);
      call5_328 <= data_out(103 downto 96);
      call6_334 <= data_out(95 downto 88);
      call7_340 <= data_out(87 downto 80);
      call8_346 <= data_out(79 downto 72);
      call9_352 <= data_out(71 downto 64);
      call22_466 <= data_out(63 downto 56);
      call25_479 <= data_out(55 downto 48);
      call30_497 <= data_out(47 downto 40);
      call36_515 <= data_out(39 downto 32);
      call42_533 <= data_out(31 downto 24);
      call48_551 <= data_out(23 downto 16);
      call54_569 <= data_out(15 downto 8);
      call60_587 <= data_out(7 downto 0);
      zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_0_gI", nreqs => 17, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 17,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_9_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_9_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_9_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_9_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_9_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_9_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_10_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_10_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_2067_start: Boolean;
  signal zeropad3D_CP_2067_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_10_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_9_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_9_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_10_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_657_call_ack_1 : boolean;
  signal LOAD_pad_660_load_0_req_1 : boolean;
  signal type_cast_1300_inst_req_0 : boolean;
  signal LOAD_pad_660_load_0_ack_1 : boolean;
  signal type_cast_1300_inst_ack_0 : boolean;
  signal LOAD_pad_660_load_0_req_0 : boolean;
  signal LOAD_out_depth_high_669_load_0_req_0 : boolean;
  signal if_stmt_1309_branch_req_0 : boolean;
  signal LOAD_out_depth_high_669_load_0_ack_0 : boolean;
  signal LOAD_depth_high_663_load_0_req_0 : boolean;
  signal LOAD_depth_high_663_load_0_ack_0 : boolean;
  signal LOAD_depth_high_663_load_0_req_1 : boolean;
  signal LOAD_depth_high_663_load_0_ack_1 : boolean;
  signal LOAD_col_high_666_load_0_ack_1 : boolean;
  signal LOAD_out_col_high_672_load_0_ack_0 : boolean;
  signal LOAD_pad_660_load_0_ack_0 : boolean;
  signal LOAD_col_high_666_load_0_req_0 : boolean;
  signal LOAD_out_col_high_672_load_0_req_0 : boolean;
  signal call_stmt_657_call_req_0 : boolean;
  signal LOAD_col_high_666_load_0_ack_0 : boolean;
  signal LOAD_out_depth_high_669_load_0_req_1 : boolean;
  signal LOAD_out_depth_high_669_load_0_ack_1 : boolean;
  signal call_stmt_657_call_req_1 : boolean;
  signal LOAD_col_high_666_load_0_req_1 : boolean;
  signal LOAD_out_col_high_672_load_0_req_1 : boolean;
  signal LOAD_out_col_high_672_load_0_ack_1 : boolean;
  signal type_cast_1218_inst_ack_0 : boolean;
  signal call_stmt_657_call_ack_0 : boolean;
  signal if_stmt_1360_branch_ack_1 : boolean;
  signal type_cast_1231_inst_ack_1 : boolean;
  signal type_cast_1300_inst_req_1 : boolean;
  signal type_cast_676_inst_req_0 : boolean;
  signal type_cast_676_inst_ack_0 : boolean;
  signal type_cast_676_inst_req_1 : boolean;
  signal type_cast_676_inst_ack_1 : boolean;
  signal type_cast_680_inst_req_0 : boolean;
  signal type_cast_680_inst_ack_0 : boolean;
  signal type_cast_680_inst_req_1 : boolean;
  signal type_cast_680_inst_ack_1 : boolean;
  signal type_cast_684_inst_req_0 : boolean;
  signal type_cast_684_inst_ack_0 : boolean;
  signal type_cast_684_inst_req_1 : boolean;
  signal type_cast_684_inst_ack_1 : boolean;
  signal type_cast_688_inst_req_0 : boolean;
  signal type_cast_688_inst_ack_0 : boolean;
  signal type_cast_688_inst_req_1 : boolean;
  signal type_cast_688_inst_ack_1 : boolean;
  signal type_cast_697_inst_req_0 : boolean;
  signal type_cast_697_inst_ack_0 : boolean;
  signal type_cast_697_inst_req_1 : boolean;
  signal type_cast_697_inst_ack_1 : boolean;
  signal type_cast_701_inst_req_0 : boolean;
  signal type_cast_701_inst_ack_0 : boolean;
  signal type_cast_701_inst_req_1 : boolean;
  signal type_cast_701_inst_ack_1 : boolean;
  signal type_cast_772_inst_req_0 : boolean;
  signal type_cast_772_inst_ack_0 : boolean;
  signal type_cast_772_inst_req_1 : boolean;
  signal type_cast_772_inst_ack_1 : boolean;
  signal if_stmt_781_branch_req_0 : boolean;
  signal if_stmt_781_branch_ack_1 : boolean;
  signal if_stmt_781_branch_ack_0 : boolean;
  signal LOAD_depth_high_1200_load_0_ack_1 : boolean;
  signal type_cast_1218_inst_req_0 : boolean;
  signal LOAD_depth_high_1200_load_0_req_1 : boolean;
  signal type_cast_1231_inst_req_1 : boolean;
  signal LOAD_row_high_789_load_0_req_0 : boolean;
  signal LOAD_row_high_789_load_0_ack_0 : boolean;
  signal LOAD_row_high_789_load_0_req_1 : boolean;
  signal LOAD_row_high_789_load_0_ack_1 : boolean;
  signal type_cast_1214_inst_ack_0 : boolean;
  signal if_stmt_1148_branch_ack_1 : boolean;
  signal type_cast_1210_inst_ack_0 : boolean;
  signal type_cast_1231_inst_ack_0 : boolean;
  signal type_cast_793_inst_req_0 : boolean;
  signal type_cast_1210_inst_req_0 : boolean;
  signal type_cast_793_inst_ack_0 : boolean;
  signal type_cast_1231_inst_req_0 : boolean;
  signal type_cast_793_inst_req_1 : boolean;
  signal type_cast_793_inst_ack_1 : boolean;
  signal if_stmt_813_branch_req_0 : boolean;
  signal if_stmt_813_branch_ack_1 : boolean;
  signal LOAD_row_high_1126_load_0_ack_1 : boolean;
  signal if_stmt_813_branch_ack_0 : boolean;
  signal type_cast_1214_inst_req_0 : boolean;
  signal type_cast_823_inst_req_0 : boolean;
  signal type_cast_823_inst_ack_0 : boolean;
  signal type_cast_823_inst_req_1 : boolean;
  signal type_cast_823_inst_ack_1 : boolean;
  signal type_cast_1300_inst_ack_1 : boolean;
  signal LOAD_row_high_1126_load_0_req_1 : boolean;
  signal LOAD_out_depth_high_1203_load_0_ack_1 : boolean;
  signal type_cast_1227_inst_ack_1 : boolean;
  signal if_stmt_832_branch_req_0 : boolean;
  signal LOAD_depth_high_1200_load_0_ack_0 : boolean;
  signal LOAD_out_depth_high_1203_load_0_req_1 : boolean;
  signal if_stmt_832_branch_ack_1 : boolean;
  signal if_stmt_832_branch_ack_0 : boolean;
  signal LOAD_depth_high_1200_load_0_req_0 : boolean;
  signal LOAD_col_high_840_load_0_req_0 : boolean;
  signal LOAD_col_high_840_load_0_ack_0 : boolean;
  signal LOAD_col_high_840_load_0_req_1 : boolean;
  signal LOAD_col_high_840_load_0_ack_1 : boolean;
  signal type_cast_1227_inst_req_1 : boolean;
  signal type_cast_844_inst_req_0 : boolean;
  signal type_cast_844_inst_ack_0 : boolean;
  signal LOAD_row_high_1126_load_0_ack_0 : boolean;
  signal type_cast_844_inst_req_1 : boolean;
  signal type_cast_844_inst_ack_1 : boolean;
  signal type_cast_1227_inst_ack_0 : boolean;
  signal if_stmt_1148_branch_req_0 : boolean;
  signal type_cast_1227_inst_req_0 : boolean;
  signal if_stmt_864_branch_req_0 : boolean;
  signal if_stmt_864_branch_ack_1 : boolean;
  signal LOAD_row_high_1126_load_0_req_0 : boolean;
  signal if_stmt_864_branch_ack_0 : boolean;
  signal LOAD_out_depth_high_1203_load_0_ack_0 : boolean;
  signal type_cast_874_inst_req_0 : boolean;
  signal type_cast_874_inst_ack_0 : boolean;
  signal LOAD_out_depth_high_1203_load_0_req_0 : boolean;
  signal type_cast_874_inst_req_1 : boolean;
  signal type_cast_874_inst_ack_1 : boolean;
  signal type_cast_1214_inst_ack_1 : boolean;
  signal type_cast_879_inst_req_0 : boolean;
  signal LOAD_out_col_high_1206_load_0_ack_1 : boolean;
  signal type_cast_879_inst_ack_0 : boolean;
  signal type_cast_879_inst_req_1 : boolean;
  signal LOAD_out_col_high_1206_load_0_req_1 : boolean;
  signal type_cast_879_inst_ack_1 : boolean;
  signal LOAD_pad_1197_load_0_ack_1 : boolean;
  signal LOAD_pad_1197_load_0_req_1 : boolean;
  signal type_cast_914_inst_req_0 : boolean;
  signal type_cast_914_inst_ack_0 : boolean;
  signal type_cast_1214_inst_req_1 : boolean;
  signal type_cast_914_inst_req_1 : boolean;
  signal type_cast_914_inst_ack_1 : boolean;
  signal type_cast_1130_inst_ack_1 : boolean;
  signal type_cast_1210_inst_ack_1 : boolean;
  signal LOAD_pad_1197_load_0_ack_0 : boolean;
  signal LOAD_pad_1197_load_0_req_0 : boolean;
  signal array_obj_ref_920_index_offset_req_0 : boolean;
  signal array_obj_ref_920_index_offset_ack_0 : boolean;
  signal type_cast_1130_inst_req_1 : boolean;
  signal array_obj_ref_920_index_offset_req_1 : boolean;
  signal array_obj_ref_920_index_offset_ack_1 : boolean;
  signal LOAD_out_col_high_1206_load_0_ack_0 : boolean;
  signal type_cast_1218_inst_ack_1 : boolean;
  signal addr_of_921_final_reg_req_0 : boolean;
  signal LOAD_out_col_high_1206_load_0_req_0 : boolean;
  signal addr_of_921_final_reg_ack_0 : boolean;
  signal type_cast_1218_inst_req_1 : boolean;
  signal addr_of_921_final_reg_req_1 : boolean;
  signal addr_of_921_final_reg_ack_1 : boolean;
  signal type_cast_1210_inst_req_1 : boolean;
  signal type_cast_1130_inst_ack_0 : boolean;
  signal type_cast_1130_inst_req_0 : boolean;
  signal type_cast_1188_inst_ack_1 : boolean;
  signal type_cast_1188_inst_req_1 : boolean;
  signal type_cast_1188_inst_ack_0 : boolean;
  signal if_stmt_1148_branch_ack_0 : boolean;
  signal ptr_deref_924_store_0_req_0 : boolean;
  signal type_cast_1188_inst_req_0 : boolean;
  signal ptr_deref_924_store_0_ack_0 : boolean;
  signal ptr_deref_924_store_0_req_1 : boolean;
  signal ptr_deref_924_store_0_ack_1 : boolean;
  signal LOAD_row_high_1831_load_0_ack_1 : boolean;
  signal type_cast_933_inst_req_0 : boolean;
  signal type_cast_933_inst_ack_0 : boolean;
  signal type_cast_1835_inst_req_1 : boolean;
  signal type_cast_933_inst_req_1 : boolean;
  signal type_cast_933_inst_ack_1 : boolean;
  signal type_cast_1835_inst_ack_1 : boolean;
  signal type_cast_997_inst_req_0 : boolean;
  signal type_cast_997_inst_ack_0 : boolean;
  signal type_cast_997_inst_req_1 : boolean;
  signal type_cast_997_inst_ack_1 : boolean;
  signal LOAD_out_col_high_1720_load_0_req_0 : boolean;
  signal type_cast_1732_inst_req_1 : boolean;
  signal type_cast_1732_inst_ack_1 : boolean;
  signal array_obj_ref_1003_index_offset_req_0 : boolean;
  signal array_obj_ref_1003_index_offset_ack_0 : boolean;
  signal array_obj_ref_1003_index_offset_req_1 : boolean;
  signal LOAD_out_col_high_1720_load_0_ack_0 : boolean;
  signal array_obj_ref_1003_index_offset_ack_1 : boolean;
  signal if_stmt_1855_branch_ack_0 : boolean;
  signal addr_of_1004_final_reg_req_0 : boolean;
  signal addr_of_1004_final_reg_ack_0 : boolean;
  signal addr_of_1004_final_reg_req_1 : boolean;
  signal addr_of_1004_final_reg_ack_1 : boolean;
  signal LOAD_out_depth_high_1717_load_0_ack_0 : boolean;
  signal if_stmt_1823_branch_req_0 : boolean;
  signal LOAD_row_high_1831_load_0_req_1 : boolean;
  signal ptr_deref_1008_load_0_req_0 : boolean;
  signal ptr_deref_1008_load_0_ack_0 : boolean;
  signal ptr_deref_1008_load_0_req_1 : boolean;
  signal ptr_deref_1008_load_0_ack_1 : boolean;
  signal type_cast_1022_inst_req_0 : boolean;
  signal type_cast_1022_inst_ack_0 : boolean;
  signal type_cast_1022_inst_req_1 : boolean;
  signal type_cast_1022_inst_ack_1 : boolean;
  signal type_cast_1741_inst_req_0 : boolean;
  signal type_cast_1741_inst_ack_0 : boolean;
  signal array_obj_ref_1028_index_offset_req_0 : boolean;
  signal array_obj_ref_1028_index_offset_ack_0 : boolean;
  signal LOAD_out_depth_high_1717_load_0_req_0 : boolean;
  signal array_obj_ref_1028_index_offset_req_1 : boolean;
  signal array_obj_ref_1028_index_offset_ack_1 : boolean;
  signal addr_of_1029_final_reg_req_0 : boolean;
  signal addr_of_1029_final_reg_ack_0 : boolean;
  signal addr_of_1029_final_reg_req_1 : boolean;
  signal addr_of_1029_final_reg_ack_1 : boolean;
  signal LOAD_row_high_1831_load_0_req_0 : boolean;
  signal LOAD_row_high_1831_load_0_ack_0 : boolean;
  signal ptr_deref_1032_store_0_req_0 : boolean;
  signal ptr_deref_1032_store_0_ack_0 : boolean;
  signal ptr_deref_1032_store_0_req_1 : boolean;
  signal ptr_deref_1032_store_0_ack_1 : boolean;
  signal type_cast_1040_inst_req_0 : boolean;
  signal type_cast_1040_inst_ack_0 : boolean;
  signal type_cast_1040_inst_req_1 : boolean;
  signal type_cast_1040_inst_ack_1 : boolean;
  signal if_stmt_1055_branch_req_0 : boolean;
  signal if_stmt_1055_branch_ack_1 : boolean;
  signal if_stmt_1055_branch_ack_0 : boolean;
  signal type_cast_1079_inst_req_0 : boolean;
  signal type_cast_1079_inst_ack_0 : boolean;
  signal type_cast_1079_inst_req_1 : boolean;
  signal type_cast_1079_inst_ack_1 : boolean;
  signal LOAD_col_high_1082_load_0_req_0 : boolean;
  signal LOAD_col_high_1082_load_0_ack_0 : boolean;
  signal LOAD_col_high_1082_load_0_req_1 : boolean;
  signal LOAD_col_high_1082_load_0_ack_1 : boolean;
  signal type_cast_1086_inst_req_0 : boolean;
  signal type_cast_1086_inst_ack_0 : boolean;
  signal type_cast_1086_inst_req_1 : boolean;
  signal type_cast_1086_inst_ack_1 : boolean;
  signal type_cast_1106_inst_req_0 : boolean;
  signal type_cast_1106_inst_ack_0 : boolean;
  signal type_cast_1106_inst_req_1 : boolean;
  signal type_cast_1106_inst_ack_1 : boolean;
  signal type_cast_1123_inst_req_0 : boolean;
  signal type_cast_1123_inst_ack_0 : boolean;
  signal type_cast_1123_inst_req_1 : boolean;
  signal type_cast_1123_inst_ack_1 : boolean;
  signal if_stmt_1309_branch_ack_1 : boolean;
  signal if_stmt_1309_branch_ack_0 : boolean;
  signal LOAD_row_high_1317_load_0_req_0 : boolean;
  signal LOAD_row_high_1317_load_0_ack_0 : boolean;
  signal LOAD_row_high_1317_load_0_req_1 : boolean;
  signal LOAD_row_high_1317_load_0_ack_1 : boolean;
  signal type_cast_1321_inst_req_0 : boolean;
  signal type_cast_1321_inst_ack_0 : boolean;
  signal type_cast_1321_inst_req_1 : boolean;
  signal type_cast_1321_inst_ack_1 : boolean;
  signal if_stmt_1341_branch_req_0 : boolean;
  signal if_stmt_1341_branch_ack_1 : boolean;
  signal if_stmt_1341_branch_ack_0 : boolean;
  signal type_cast_1351_inst_req_0 : boolean;
  signal type_cast_1351_inst_ack_0 : boolean;
  signal type_cast_1351_inst_req_1 : boolean;
  signal type_cast_1351_inst_ack_1 : boolean;
  signal if_stmt_1360_branch_req_0 : boolean;
  signal type_cast_3813_inst_ack_0 : boolean;
  signal if_stmt_1360_branch_ack_0 : boolean;
  signal LOAD_col_high_1368_load_0_req_0 : boolean;
  signal LOAD_col_high_1368_load_0_ack_0 : boolean;
  signal LOAD_col_high_1368_load_0_req_1 : boolean;
  signal LOAD_col_high_1368_load_0_ack_1 : boolean;
  signal type_cast_1372_inst_req_0 : boolean;
  signal type_cast_1372_inst_ack_0 : boolean;
  signal type_cast_1372_inst_req_1 : boolean;
  signal type_cast_1372_inst_ack_1 : boolean;
  signal if_stmt_1386_branch_req_0 : boolean;
  signal if_stmt_1386_branch_ack_1 : boolean;
  signal if_stmt_1386_branch_ack_0 : boolean;
  signal type_cast_1835_inst_ack_0 : boolean;
  signal type_cast_1396_inst_req_0 : boolean;
  signal type_cast_1814_inst_ack_1 : boolean;
  signal type_cast_1396_inst_ack_0 : boolean;
  signal type_cast_1741_inst_ack_1 : boolean;
  signal type_cast_1835_inst_req_0 : boolean;
  signal type_cast_1396_inst_req_1 : boolean;
  signal type_cast_1814_inst_req_1 : boolean;
  signal type_cast_1396_inst_ack_1 : boolean;
  signal type_cast_1732_inst_ack_0 : boolean;
  signal type_cast_1732_inst_req_0 : boolean;
  signal type_cast_1401_inst_req_0 : boolean;
  signal type_cast_1401_inst_ack_0 : boolean;
  signal type_cast_1401_inst_req_1 : boolean;
  signal type_cast_1401_inst_ack_1 : boolean;
  signal type_cast_1814_inst_ack_0 : boolean;
  signal type_cast_1435_inst_req_0 : boolean;
  signal type_cast_1814_inst_req_0 : boolean;
  signal type_cast_1435_inst_ack_0 : boolean;
  signal type_cast_1435_inst_req_1 : boolean;
  signal type_cast_1435_inst_ack_1 : boolean;
  signal type_cast_1728_inst_ack_1 : boolean;
  signal type_cast_1728_inst_req_1 : boolean;
  signal array_obj_ref_1441_index_offset_req_0 : boolean;
  signal array_obj_ref_1441_index_offset_ack_0 : boolean;
  signal array_obj_ref_1441_index_offset_req_1 : boolean;
  signal array_obj_ref_1441_index_offset_ack_1 : boolean;
  signal if_stmt_1855_branch_ack_1 : boolean;
  signal type_cast_1728_inst_ack_0 : boolean;
  signal addr_of_1442_final_reg_req_0 : boolean;
  signal addr_of_1442_final_reg_ack_0 : boolean;
  signal addr_of_1442_final_reg_req_1 : boolean;
  signal addr_of_1442_final_reg_ack_1 : boolean;
  signal if_stmt_1823_branch_ack_0 : boolean;
  signal type_cast_1728_inst_req_0 : boolean;
  signal type_cast_1724_inst_ack_1 : boolean;
  signal type_cast_1724_inst_req_1 : boolean;
  signal type_cast_1745_inst_ack_1 : boolean;
  signal type_cast_1724_inst_ack_0 : boolean;
  signal type_cast_1745_inst_req_1 : boolean;
  signal LOAD_out_col_high_1720_load_0_ack_1 : boolean;
  signal ptr_deref_1445_store_0_req_0 : boolean;
  signal type_cast_1724_inst_req_0 : boolean;
  signal ptr_deref_1445_store_0_ack_0 : boolean;
  signal LOAD_out_col_high_1720_load_0_req_1 : boolean;
  signal ptr_deref_1445_store_0_req_1 : boolean;
  signal ptr_deref_1445_store_0_ack_1 : boolean;
  signal if_stmt_1855_branch_req_0 : boolean;
  signal type_cast_1745_inst_ack_0 : boolean;
  signal type_cast_1454_inst_req_0 : boolean;
  signal type_cast_1745_inst_req_0 : boolean;
  signal type_cast_1454_inst_ack_0 : boolean;
  signal type_cast_1741_inst_req_1 : boolean;
  signal type_cast_1454_inst_req_1 : boolean;
  signal type_cast_1454_inst_ack_1 : boolean;
  signal LOAD_out_depth_high_1717_load_0_ack_1 : boolean;
  signal LOAD_out_depth_high_1717_load_0_req_1 : boolean;
  signal if_stmt_1823_branch_ack_1 : boolean;
  signal type_cast_1518_inst_req_0 : boolean;
  signal type_cast_1518_inst_ack_0 : boolean;
  signal type_cast_1518_inst_req_1 : boolean;
  signal type_cast_1518_inst_ack_1 : boolean;
  signal type_cast_2375_inst_req_0 : boolean;
  signal array_obj_ref_1524_index_offset_req_0 : boolean;
  signal array_obj_ref_1524_index_offset_ack_0 : boolean;
  signal array_obj_ref_1524_index_offset_req_1 : boolean;
  signal array_obj_ref_1524_index_offset_ack_1 : boolean;
  signal type_cast_2375_inst_ack_0 : boolean;
  signal addr_of_1525_final_reg_req_0 : boolean;
  signal addr_of_1525_final_reg_ack_0 : boolean;
  signal addr_of_1525_final_reg_req_1 : boolean;
  signal addr_of_1525_final_reg_ack_1 : boolean;
  signal type_cast_2426_inst_ack_0 : boolean;
  signal type_cast_2282_inst_req_1 : boolean;
  signal type_cast_2375_inst_req_1 : boolean;
  signal type_cast_2375_inst_ack_1 : boolean;
  signal if_stmt_2414_branch_ack_1 : boolean;
  signal ptr_deref_1529_load_0_req_0 : boolean;
  signal ptr_deref_1529_load_0_ack_0 : boolean;
  signal ptr_deref_1529_load_0_req_1 : boolean;
  signal ptr_deref_1529_load_0_ack_1 : boolean;
  signal type_cast_2282_inst_ack_1 : boolean;
  signal type_cast_1543_inst_req_0 : boolean;
  signal type_cast_1543_inst_ack_0 : boolean;
  signal type_cast_1543_inst_req_1 : boolean;
  signal type_cast_1543_inst_ack_1 : boolean;
  signal if_stmt_2363_branch_req_0 : boolean;
  signal array_obj_ref_1549_index_offset_req_0 : boolean;
  signal array_obj_ref_1549_index_offset_ack_0 : boolean;
  signal if_stmt_2395_branch_req_0 : boolean;
  signal array_obj_ref_1549_index_offset_req_1 : boolean;
  signal array_obj_ref_1549_index_offset_ack_1 : boolean;
  signal if_stmt_2414_branch_ack_0 : boolean;
  signal addr_of_1550_final_reg_req_0 : boolean;
  signal addr_of_1550_final_reg_ack_0 : boolean;
  signal addr_of_1550_final_reg_req_1 : boolean;
  signal addr_of_1550_final_reg_ack_1 : boolean;
  signal type_cast_2426_inst_req_1 : boolean;
  signal type_cast_2426_inst_ack_1 : boolean;
  signal if_stmt_2395_branch_ack_1 : boolean;
  signal ptr_deref_1553_store_0_req_0 : boolean;
  signal ptr_deref_1553_store_0_ack_0 : boolean;
  signal if_stmt_2363_branch_ack_1 : boolean;
  signal ptr_deref_1553_store_0_req_1 : boolean;
  signal if_stmt_2395_branch_ack_0 : boolean;
  signal ptr_deref_1553_store_0_ack_1 : boolean;
  signal type_cast_2426_inst_req_0 : boolean;
  signal type_cast_1561_inst_req_0 : boolean;
  signal type_cast_1561_inst_ack_0 : boolean;
  signal type_cast_1561_inst_req_1 : boolean;
  signal type_cast_1561_inst_ack_1 : boolean;
  signal if_stmt_2363_branch_ack_0 : boolean;
  signal type_cast_2405_inst_req_0 : boolean;
  signal LOAD_col_high_2422_load_0_req_0 : boolean;
  signal if_stmt_1576_branch_req_0 : boolean;
  signal if_stmt_1576_branch_ack_1 : boolean;
  signal type_cast_2286_inst_req_0 : boolean;
  signal if_stmt_1576_branch_ack_0 : boolean;
  signal type_cast_2405_inst_ack_0 : boolean;
  signal type_cast_2286_inst_ack_0 : boolean;
  signal type_cast_1600_inst_req_0 : boolean;
  signal type_cast_1600_inst_ack_0 : boolean;
  signal type_cast_1600_inst_req_1 : boolean;
  signal type_cast_1600_inst_ack_1 : boolean;
  signal LOAD_col_high_1603_load_0_req_0 : boolean;
  signal LOAD_col_high_1603_load_0_ack_0 : boolean;
  signal LOAD_col_high_1603_load_0_req_1 : boolean;
  signal LOAD_col_high_1603_load_0_ack_1 : boolean;
  signal type_cast_1607_inst_req_0 : boolean;
  signal type_cast_1607_inst_ack_0 : boolean;
  signal type_cast_1607_inst_req_1 : boolean;
  signal type_cast_1607_inst_ack_1 : boolean;
  signal type_cast_1621_inst_req_0 : boolean;
  signal type_cast_1621_inst_ack_0 : boolean;
  signal type_cast_1621_inst_req_1 : boolean;
  signal type_cast_1621_inst_ack_1 : boolean;
  signal type_cast_1637_inst_req_0 : boolean;
  signal type_cast_1637_inst_ack_0 : boolean;
  signal type_cast_1637_inst_req_1 : boolean;
  signal type_cast_1637_inst_ack_1 : boolean;
  signal LOAD_row_high_1640_load_0_req_0 : boolean;
  signal LOAD_row_high_1640_load_0_ack_0 : boolean;
  signal LOAD_row_high_1640_load_0_req_1 : boolean;
  signal LOAD_row_high_1640_load_0_ack_1 : boolean;
  signal type_cast_1644_inst_req_0 : boolean;
  signal type_cast_1644_inst_ack_0 : boolean;
  signal type_cast_1644_inst_req_1 : boolean;
  signal type_cast_1644_inst_ack_1 : boolean;
  signal if_stmt_1662_branch_req_0 : boolean;
  signal if_stmt_1662_branch_ack_1 : boolean;
  signal if_stmt_1662_branch_ack_0 : boolean;
  signal type_cast_1702_inst_req_0 : boolean;
  signal type_cast_1702_inst_ack_0 : boolean;
  signal type_cast_1702_inst_req_1 : boolean;
  signal type_cast_1702_inst_ack_1 : boolean;
  signal LOAD_pad_1711_load_0_req_0 : boolean;
  signal LOAD_pad_1711_load_0_ack_0 : boolean;
  signal LOAD_pad_1711_load_0_req_1 : boolean;
  signal LOAD_pad_1711_load_0_ack_1 : boolean;
  signal LOAD_depth_high_1714_load_0_req_0 : boolean;
  signal LOAD_depth_high_1714_load_0_ack_0 : boolean;
  signal LOAD_depth_high_1714_load_0_req_1 : boolean;
  signal LOAD_depth_high_1714_load_0_ack_1 : boolean;
  signal type_cast_1865_inst_req_0 : boolean;
  signal type_cast_1865_inst_ack_0 : boolean;
  signal type_cast_1865_inst_req_1 : boolean;
  signal type_cast_1865_inst_ack_1 : boolean;
  signal if_stmt_1874_branch_req_0 : boolean;
  signal if_stmt_1874_branch_ack_1 : boolean;
  signal if_stmt_1874_branch_ack_0 : boolean;
  signal LOAD_col_high_1882_load_0_req_0 : boolean;
  signal LOAD_col_high_1882_load_0_ack_0 : boolean;
  signal LOAD_col_high_1882_load_0_req_1 : boolean;
  signal LOAD_col_high_1882_load_0_ack_1 : boolean;
  signal type_cast_1886_inst_req_0 : boolean;
  signal type_cast_1886_inst_ack_0 : boolean;
  signal type_cast_1886_inst_req_1 : boolean;
  signal type_cast_1886_inst_ack_1 : boolean;
  signal if_stmt_1906_branch_req_0 : boolean;
  signal if_stmt_1906_branch_ack_1 : boolean;
  signal if_stmt_1906_branch_ack_0 : boolean;
  signal type_cast_1916_inst_req_0 : boolean;
  signal type_cast_1916_inst_ack_0 : boolean;
  signal type_cast_1916_inst_req_1 : boolean;
  signal type_cast_1916_inst_ack_1 : boolean;
  signal type_cast_1921_inst_req_0 : boolean;
  signal type_cast_1921_inst_ack_0 : boolean;
  signal type_cast_1921_inst_req_1 : boolean;
  signal type_cast_1921_inst_ack_1 : boolean;
  signal type_cast_1955_inst_req_0 : boolean;
  signal type_cast_1955_inst_ack_0 : boolean;
  signal type_cast_1955_inst_req_1 : boolean;
  signal type_cast_1955_inst_ack_1 : boolean;
  signal array_obj_ref_1961_index_offset_req_0 : boolean;
  signal array_obj_ref_1961_index_offset_ack_0 : boolean;
  signal array_obj_ref_1961_index_offset_req_1 : boolean;
  signal array_obj_ref_1961_index_offset_ack_1 : boolean;
  signal addr_of_1962_final_reg_req_0 : boolean;
  signal addr_of_1962_final_reg_ack_0 : boolean;
  signal addr_of_1962_final_reg_req_1 : boolean;
  signal addr_of_1962_final_reg_ack_1 : boolean;
  signal if_stmt_2414_branch_req_0 : boolean;
  signal LOAD_col_high_2422_load_0_ack_1 : boolean;
  signal ptr_deref_1965_store_0_req_0 : boolean;
  signal ptr_deref_1965_store_0_ack_0 : boolean;
  signal type_cast_2282_inst_ack_0 : boolean;
  signal ptr_deref_1965_store_0_req_1 : boolean;
  signal ptr_deref_1965_store_0_ack_1 : boolean;
  signal type_cast_2354_inst_ack_1 : boolean;
  signal type_cast_2354_inst_req_1 : boolean;
  signal type_cast_2282_inst_req_0 : boolean;
  signal LOAD_row_high_2371_load_0_ack_1 : boolean;
  signal LOAD_row_high_2371_load_0_req_1 : boolean;
  signal type_cast_1974_inst_req_0 : boolean;
  signal type_cast_1974_inst_ack_0 : boolean;
  signal type_cast_1974_inst_req_1 : boolean;
  signal type_cast_1974_inst_ack_1 : boolean;
  signal type_cast_2286_inst_ack_1 : boolean;
  signal type_cast_2286_inst_req_1 : boolean;
  signal LOAD_col_high_2422_load_0_req_1 : boolean;
  signal type_cast_2038_inst_req_0 : boolean;
  signal type_cast_2038_inst_ack_0 : boolean;
  signal type_cast_2038_inst_req_1 : boolean;
  signal type_cast_2405_inst_ack_1 : boolean;
  signal type_cast_2038_inst_ack_1 : boolean;
  signal LOAD_row_high_2371_load_0_ack_0 : boolean;
  signal LOAD_row_high_2371_load_0_req_0 : boolean;
  signal array_obj_ref_2044_index_offset_req_0 : boolean;
  signal type_cast_2405_inst_req_1 : boolean;
  signal array_obj_ref_2044_index_offset_ack_0 : boolean;
  signal type_cast_2354_inst_ack_0 : boolean;
  signal array_obj_ref_2044_index_offset_req_1 : boolean;
  signal array_obj_ref_2044_index_offset_ack_1 : boolean;
  signal LOAD_col_high_2422_load_0_ack_0 : boolean;
  signal type_cast_2354_inst_req_0 : boolean;
  signal addr_of_2045_final_reg_req_0 : boolean;
  signal addr_of_2045_final_reg_ack_0 : boolean;
  signal addr_of_2045_final_reg_req_1 : boolean;
  signal addr_of_2045_final_reg_ack_1 : boolean;
  signal LOAD_pad_2765_load_0_ack_1 : boolean;
  signal if_stmt_2934_branch_ack_0 : boolean;
  signal type_cast_2786_inst_req_1 : boolean;
  signal type_cast_2786_inst_ack_1 : boolean;
  signal ptr_deref_2049_load_0_req_0 : boolean;
  signal ptr_deref_2049_load_0_ack_0 : boolean;
  signal ptr_deref_2049_load_0_req_1 : boolean;
  signal ptr_deref_2049_load_0_ack_1 : boolean;
  signal type_cast_2063_inst_req_0 : boolean;
  signal LOAD_out_depth_high_2771_load_0_req_1 : boolean;
  signal type_cast_2063_inst_ack_0 : boolean;
  signal if_stmt_2966_branch_ack_0 : boolean;
  signal type_cast_2063_inst_req_1 : boolean;
  signal type_cast_2063_inst_ack_1 : boolean;
  signal LOAD_out_depth_high_2771_load_0_ack_1 : boolean;
  signal type_cast_2795_inst_req_0 : boolean;
  signal array_obj_ref_2069_index_offset_req_0 : boolean;
  signal array_obj_ref_2069_index_offset_ack_0 : boolean;
  signal array_obj_ref_2069_index_offset_req_1 : boolean;
  signal type_cast_2795_inst_ack_0 : boolean;
  signal array_obj_ref_2069_index_offset_ack_1 : boolean;
  signal addr_of_2070_final_reg_req_0 : boolean;
  signal addr_of_2070_final_reg_ack_0 : boolean;
  signal addr_of_2070_final_reg_req_1 : boolean;
  signal addr_of_2070_final_reg_ack_1 : boolean;
  signal type_cast_2795_inst_req_1 : boolean;
  signal type_cast_2795_inst_ack_1 : boolean;
  signal type_cast_2889_inst_req_0 : boolean;
  signal ptr_deref_2073_store_0_req_0 : boolean;
  signal ptr_deref_2073_store_0_ack_0 : boolean;
  signal LOAD_col_high_2942_load_0_req_0 : boolean;
  signal ptr_deref_2073_store_0_req_1 : boolean;
  signal ptr_deref_2073_store_0_ack_1 : boolean;
  signal LOAD_out_col_high_2774_load_0_req_1 : boolean;
  signal type_cast_2081_inst_req_0 : boolean;
  signal type_cast_2889_inst_ack_0 : boolean;
  signal type_cast_2081_inst_ack_0 : boolean;
  signal type_cast_2081_inst_req_1 : boolean;
  signal type_cast_2081_inst_ack_1 : boolean;
  signal if_stmt_2877_branch_req_0 : boolean;
  signal LOAD_out_depth_high_2771_load_0_req_0 : boolean;
  signal if_stmt_2096_branch_req_0 : boolean;
  signal if_stmt_2096_branch_ack_1 : boolean;
  signal LOAD_out_depth_high_2771_load_0_ack_0 : boolean;
  signal if_stmt_2096_branch_ack_0 : boolean;
  signal LOAD_out_col_high_2774_load_0_ack_1 : boolean;
  signal type_cast_2120_inst_req_0 : boolean;
  signal type_cast_2120_inst_ack_0 : boolean;
  signal type_cast_2120_inst_req_1 : boolean;
  signal type_cast_2120_inst_ack_1 : boolean;
  signal type_cast_2799_inst_req_0 : boolean;
  signal type_cast_2799_inst_ack_0 : boolean;
  signal LOAD_col_high_2123_load_0_req_0 : boolean;
  signal LOAD_col_high_2123_load_0_ack_0 : boolean;
  signal LOAD_col_high_2123_load_0_req_1 : boolean;
  signal LOAD_col_high_2123_load_0_ack_1 : boolean;
  signal LOAD_col_high_2942_load_0_ack_0 : boolean;
  signal type_cast_2127_inst_req_0 : boolean;
  signal type_cast_2127_inst_ack_0 : boolean;
  signal type_cast_2127_inst_req_1 : boolean;
  signal type_cast_2127_inst_ack_1 : boolean;
  signal type_cast_3015_inst_ack_1 : boolean;
  signal type_cast_2147_inst_req_0 : boolean;
  signal type_cast_2147_inst_ack_0 : boolean;
  signal type_cast_2147_inst_req_1 : boolean;
  signal type_cast_2889_inst_req_1 : boolean;
  signal type_cast_2147_inst_ack_1 : boolean;
  signal type_cast_2889_inst_ack_1 : boolean;
  signal type_cast_2799_inst_req_1 : boolean;
  signal type_cast_2799_inst_ack_1 : boolean;
  signal type_cast_2164_inst_req_0 : boolean;
  signal type_cast_2164_inst_ack_0 : boolean;
  signal type_cast_2164_inst_req_1 : boolean;
  signal type_cast_2164_inst_ack_1 : boolean;
  signal LOAD_row_high_2167_load_0_req_0 : boolean;
  signal LOAD_row_high_2167_load_0_ack_0 : boolean;
  signal LOAD_row_high_2167_load_0_req_1 : boolean;
  signal LOAD_row_high_2167_load_0_ack_1 : boolean;
  signal type_cast_2171_inst_req_0 : boolean;
  signal type_cast_2171_inst_ack_0 : boolean;
  signal type_cast_2171_inst_req_1 : boolean;
  signal type_cast_2171_inst_ack_1 : boolean;
  signal if_stmt_2189_branch_req_0 : boolean;
  signal if_stmt_2189_branch_ack_1 : boolean;
  signal if_stmt_2189_branch_ack_0 : boolean;
  signal type_cast_2233_inst_req_0 : boolean;
  signal type_cast_2233_inst_ack_0 : boolean;
  signal type_cast_2233_inst_req_1 : boolean;
  signal type_cast_2233_inst_ack_1 : boolean;
  signal type_cast_2243_inst_req_0 : boolean;
  signal type_cast_2243_inst_ack_0 : boolean;
  signal type_cast_2243_inst_req_1 : boolean;
  signal type_cast_2243_inst_ack_1 : boolean;
  signal LOAD_pad_2252_load_0_req_0 : boolean;
  signal LOAD_pad_2252_load_0_ack_0 : boolean;
  signal LOAD_pad_2252_load_0_req_1 : boolean;
  signal LOAD_pad_2252_load_0_ack_1 : boolean;
  signal LOAD_depth_high_2255_load_0_req_0 : boolean;
  signal LOAD_depth_high_2255_load_0_ack_0 : boolean;
  signal LOAD_depth_high_2255_load_0_req_1 : boolean;
  signal LOAD_depth_high_2255_load_0_ack_1 : boolean;
  signal LOAD_out_depth_high_2258_load_0_req_0 : boolean;
  signal LOAD_out_depth_high_2258_load_0_ack_0 : boolean;
  signal LOAD_out_depth_high_2258_load_0_req_1 : boolean;
  signal LOAD_out_depth_high_2258_load_0_ack_1 : boolean;
  signal LOAD_out_col_high_2261_load_0_req_0 : boolean;
  signal LOAD_out_col_high_2261_load_0_ack_0 : boolean;
  signal LOAD_out_col_high_2261_load_0_req_1 : boolean;
  signal LOAD_out_col_high_2261_load_0_ack_1 : boolean;
  signal type_cast_2265_inst_req_0 : boolean;
  signal type_cast_2265_inst_ack_0 : boolean;
  signal type_cast_2265_inst_req_1 : boolean;
  signal type_cast_2265_inst_ack_1 : boolean;
  signal type_cast_2269_inst_req_0 : boolean;
  signal type_cast_2269_inst_ack_0 : boolean;
  signal type_cast_2269_inst_req_1 : boolean;
  signal type_cast_2269_inst_ack_1 : boolean;
  signal type_cast_2273_inst_req_0 : boolean;
  signal type_cast_2273_inst_ack_0 : boolean;
  signal type_cast_2273_inst_req_1 : boolean;
  signal type_cast_2273_inst_ack_1 : boolean;
  signal if_stmt_2440_branch_req_0 : boolean;
  signal if_stmt_2440_branch_ack_1 : boolean;
  signal if_stmt_2440_branch_ack_0 : boolean;
  signal type_cast_2450_inst_req_0 : boolean;
  signal type_cast_2450_inst_ack_0 : boolean;
  signal type_cast_2450_inst_req_1 : boolean;
  signal type_cast_2450_inst_ack_1 : boolean;
  signal type_cast_2455_inst_req_0 : boolean;
  signal type_cast_2455_inst_ack_0 : boolean;
  signal type_cast_2455_inst_req_1 : boolean;
  signal type_cast_2455_inst_ack_1 : boolean;
  signal type_cast_2489_inst_req_0 : boolean;
  signal type_cast_2489_inst_ack_0 : boolean;
  signal type_cast_2489_inst_req_1 : boolean;
  signal type_cast_2489_inst_ack_1 : boolean;
  signal array_obj_ref_2495_index_offset_req_0 : boolean;
  signal array_obj_ref_2495_index_offset_ack_0 : boolean;
  signal array_obj_ref_2495_index_offset_req_1 : boolean;
  signal array_obj_ref_2495_index_offset_ack_1 : boolean;
  signal addr_of_2496_final_reg_req_0 : boolean;
  signal addr_of_2496_final_reg_ack_0 : boolean;
  signal addr_of_2496_final_reg_req_1 : boolean;
  signal addr_of_2496_final_reg_ack_1 : boolean;
  signal ptr_deref_2499_store_0_req_0 : boolean;
  signal ptr_deref_2499_store_0_ack_0 : boolean;
  signal ptr_deref_2499_store_0_req_1 : boolean;
  signal ptr_deref_2499_store_0_ack_1 : boolean;
  signal type_cast_2508_inst_req_0 : boolean;
  signal type_cast_2508_inst_ack_0 : boolean;
  signal type_cast_2508_inst_req_1 : boolean;
  signal type_cast_2508_inst_ack_1 : boolean;
  signal type_cast_2572_inst_req_0 : boolean;
  signal type_cast_2572_inst_ack_0 : boolean;
  signal type_cast_2572_inst_req_1 : boolean;
  signal type_cast_2572_inst_ack_1 : boolean;
  signal array_obj_ref_2578_index_offset_req_0 : boolean;
  signal array_obj_ref_2578_index_offset_ack_0 : boolean;
  signal array_obj_ref_2578_index_offset_req_1 : boolean;
  signal array_obj_ref_2578_index_offset_ack_1 : boolean;
  signal addr_of_2579_final_reg_req_0 : boolean;
  signal addr_of_2579_final_reg_ack_0 : boolean;
  signal if_stmt_2966_branch_ack_1 : boolean;
  signal addr_of_2579_final_reg_req_1 : boolean;
  signal addr_of_2579_final_reg_ack_1 : boolean;
  signal type_cast_3015_inst_req_1 : boolean;
  signal if_stmt_2934_branch_ack_1 : boolean;
  signal if_stmt_2934_branch_req_0 : boolean;
  signal type_cast_2868_inst_ack_1 : boolean;
  signal LOAD_row_high_2885_load_0_ack_1 : boolean;
  signal ptr_deref_2583_load_0_req_0 : boolean;
  signal ptr_deref_2583_load_0_ack_0 : boolean;
  signal LOAD_row_high_2885_load_0_req_1 : boolean;
  signal ptr_deref_2583_load_0_req_1 : boolean;
  signal ptr_deref_2583_load_0_ack_1 : boolean;
  signal LOAD_depth_high_2768_load_0_ack_1 : boolean;
  signal LOAD_depth_high_2768_load_0_req_1 : boolean;
  signal LOAD_pad_2765_load_0_req_1 : boolean;
  signal type_cast_2597_inst_req_0 : boolean;
  signal type_cast_2597_inst_ack_0 : boolean;
  signal type_cast_2868_inst_req_1 : boolean;
  signal if_stmt_2966_branch_req_0 : boolean;
  signal type_cast_2597_inst_req_1 : boolean;
  signal type_cast_2597_inst_ack_1 : boolean;
  signal type_cast_3015_inst_ack_0 : boolean;
  signal type_cast_3015_inst_req_0 : boolean;
  signal type_cast_2925_inst_ack_1 : boolean;
  signal type_cast_2925_inst_req_1 : boolean;
  signal type_cast_2786_inst_ack_0 : boolean;
  signal type_cast_2925_inst_ack_0 : boolean;
  signal type_cast_2786_inst_req_0 : boolean;
  signal array_obj_ref_2603_index_offset_req_0 : boolean;
  signal array_obj_ref_2603_index_offset_ack_0 : boolean;
  signal array_obj_ref_2603_index_offset_req_1 : boolean;
  signal array_obj_ref_2603_index_offset_ack_1 : boolean;
  signal type_cast_2976_inst_ack_1 : boolean;
  signal type_cast_2976_inst_req_1 : boolean;
  signal LOAD_row_high_2885_load_0_ack_0 : boolean;
  signal addr_of_2604_final_reg_req_0 : boolean;
  signal addr_of_2604_final_reg_ack_0 : boolean;
  signal LOAD_row_high_2885_load_0_req_0 : boolean;
  signal addr_of_2604_final_reg_req_1 : boolean;
  signal addr_of_2604_final_reg_ack_1 : boolean;
  signal type_cast_2925_inst_req_0 : boolean;
  signal type_cast_2782_inst_ack_1 : boolean;
  signal type_cast_2782_inst_req_1 : boolean;
  signal type_cast_2868_inst_ack_0 : boolean;
  signal ptr_deref_2607_store_0_req_0 : boolean;
  signal ptr_deref_2607_store_0_ack_0 : boolean;
  signal LOAD_depth_high_2768_load_0_ack_0 : boolean;
  signal ptr_deref_2607_store_0_req_1 : boolean;
  signal ptr_deref_2607_store_0_ack_1 : boolean;
  signal LOAD_depth_high_2768_load_0_req_0 : boolean;
  signal type_cast_2615_inst_req_0 : boolean;
  signal type_cast_2615_inst_ack_0 : boolean;
  signal type_cast_2868_inst_req_0 : boolean;
  signal type_cast_2615_inst_req_1 : boolean;
  signal type_cast_2615_inst_ack_1 : boolean;
  signal type_cast_2946_inst_ack_1 : boolean;
  signal type_cast_2946_inst_req_1 : boolean;
  signal if_stmt_2630_branch_req_0 : boolean;
  signal type_cast_2976_inst_ack_0 : boolean;
  signal type_cast_2782_inst_ack_0 : boolean;
  signal if_stmt_2630_branch_ack_1 : boolean;
  signal if_stmt_2630_branch_ack_0 : boolean;
  signal LOAD_out_col_high_2774_load_0_ack_0 : boolean;
  signal if_stmt_2915_branch_ack_0 : boolean;
  signal LOAD_out_col_high_2774_load_0_req_0 : boolean;
  signal type_cast_2654_inst_req_0 : boolean;
  signal type_cast_2654_inst_ack_0 : boolean;
  signal type_cast_2946_inst_ack_0 : boolean;
  signal type_cast_2946_inst_req_0 : boolean;
  signal type_cast_2654_inst_req_1 : boolean;
  signal type_cast_2654_inst_ack_1 : boolean;
  signal type_cast_2981_inst_ack_1 : boolean;
  signal if_stmt_2915_branch_ack_1 : boolean;
  signal type_cast_2782_inst_req_0 : boolean;
  signal LOAD_col_high_2657_load_0_req_0 : boolean;
  signal LOAD_col_high_2657_load_0_ack_0 : boolean;
  signal LOAD_col_high_2657_load_0_req_1 : boolean;
  signal LOAD_col_high_2657_load_0_ack_1 : boolean;
  signal type_cast_2778_inst_ack_1 : boolean;
  signal type_cast_2976_inst_req_0 : boolean;
  signal type_cast_2778_inst_req_1 : boolean;
  signal type_cast_2661_inst_req_0 : boolean;
  signal type_cast_2661_inst_ack_0 : boolean;
  signal type_cast_2661_inst_req_1 : boolean;
  signal type_cast_2661_inst_ack_1 : boolean;
  signal type_cast_2981_inst_req_1 : boolean;
  signal if_stmt_2915_branch_req_0 : boolean;
  signal type_cast_2675_inst_req_0 : boolean;
  signal type_cast_2675_inst_ack_0 : boolean;
  signal type_cast_2675_inst_req_1 : boolean;
  signal type_cast_2675_inst_ack_1 : boolean;
  signal type_cast_2981_inst_ack_0 : boolean;
  signal if_stmt_2877_branch_ack_0 : boolean;
  signal type_cast_2691_inst_req_0 : boolean;
  signal type_cast_2691_inst_ack_0 : boolean;
  signal LOAD_col_high_2942_load_0_ack_1 : boolean;
  signal type_cast_2691_inst_req_1 : boolean;
  signal type_cast_2691_inst_ack_1 : boolean;
  signal type_cast_2981_inst_req_0 : boolean;
  signal type_cast_2778_inst_ack_0 : boolean;
  signal LOAD_col_high_2942_load_0_req_1 : boolean;
  signal LOAD_row_high_2694_load_0_req_0 : boolean;
  signal type_cast_2778_inst_req_0 : boolean;
  signal LOAD_row_high_2694_load_0_ack_0 : boolean;
  signal LOAD_row_high_2694_load_0_req_1 : boolean;
  signal LOAD_row_high_2694_load_0_ack_1 : boolean;
  signal if_stmt_2877_branch_ack_1 : boolean;
  signal type_cast_2698_inst_req_0 : boolean;
  signal type_cast_2698_inst_ack_0 : boolean;
  signal type_cast_2698_inst_req_1 : boolean;
  signal type_cast_2698_inst_ack_1 : boolean;
  signal LOAD_col_high_3494_load_0_req_0 : boolean;
  signal type_cast_3352_inst_req_1 : boolean;
  signal if_stmt_2716_branch_req_0 : boolean;
  signal type_cast_3339_inst_req_1 : boolean;
  signal type_cast_3352_inst_ack_1 : boolean;
  signal type_cast_3339_inst_ack_1 : boolean;
  signal if_stmt_2716_branch_ack_1 : boolean;
  signal if_stmt_2716_branch_ack_0 : boolean;
  signal if_stmt_3467_branch_ack_1 : boolean;
  signal type_cast_2756_inst_req_0 : boolean;
  signal type_cast_2756_inst_ack_0 : boolean;
  signal type_cast_2756_inst_req_1 : boolean;
  signal type_cast_2756_inst_ack_1 : boolean;
  signal LOAD_pad_2765_load_0_req_0 : boolean;
  signal LOAD_pad_2765_load_0_ack_0 : boolean;
  signal array_obj_ref_3021_index_offset_req_0 : boolean;
  signal array_obj_ref_3021_index_offset_ack_0 : boolean;
  signal array_obj_ref_3021_index_offset_req_1 : boolean;
  signal array_obj_ref_3021_index_offset_ack_1 : boolean;
  signal addr_of_3022_final_reg_req_0 : boolean;
  signal addr_of_3022_final_reg_ack_0 : boolean;
  signal addr_of_3022_final_reg_req_1 : boolean;
  signal addr_of_3022_final_reg_ack_1 : boolean;
  signal ptr_deref_3025_store_0_req_0 : boolean;
  signal ptr_deref_3025_store_0_ack_0 : boolean;
  signal ptr_deref_3025_store_0_req_1 : boolean;
  signal ptr_deref_3025_store_0_ack_1 : boolean;
  signal type_cast_3034_inst_req_0 : boolean;
  signal type_cast_3034_inst_ack_0 : boolean;
  signal type_cast_3034_inst_req_1 : boolean;
  signal type_cast_3034_inst_ack_1 : boolean;
  signal type_cast_3098_inst_req_0 : boolean;
  signal type_cast_3098_inst_ack_0 : boolean;
  signal type_cast_3098_inst_req_1 : boolean;
  signal type_cast_3098_inst_ack_1 : boolean;
  signal type_cast_4048_inst_ack_0 : boolean;
  signal if_stmt_3512_branch_ack_0 : boolean;
  signal if_stmt_3467_branch_req_0 : boolean;
  signal LOAD_row_high_3437_load_0_ack_0 : boolean;
  signal array_obj_ref_3567_index_offset_req_1 : boolean;
  signal LOAD_row_high_3437_load_0_req_0 : boolean;
  signal array_obj_ref_3104_index_offset_req_0 : boolean;
  signal array_obj_ref_3104_index_offset_ack_0 : boolean;
  signal array_obj_ref_3104_index_offset_req_1 : boolean;
  signal array_obj_ref_3104_index_offset_ack_1 : boolean;
  signal type_cast_3522_inst_ack_1 : boolean;
  signal type_cast_3348_inst_ack_0 : boolean;
  signal array_obj_ref_3567_index_offset_ack_0 : boolean;
  signal addr_of_3105_final_reg_req_0 : boolean;
  signal addr_of_3105_final_reg_ack_0 : boolean;
  signal addr_of_3105_final_reg_req_1 : boolean;
  signal addr_of_3105_final_reg_ack_1 : boolean;
  signal if_stmt_3512_branch_ack_1 : boolean;
  signal type_cast_3339_inst_ack_0 : boolean;
  signal type_cast_3339_inst_req_0 : boolean;
  signal ptr_deref_3109_load_0_req_0 : boolean;
  signal ptr_deref_3109_load_0_ack_0 : boolean;
  signal type_cast_3352_inst_ack_0 : boolean;
  signal ptr_deref_3109_load_0_req_1 : boolean;
  signal ptr_deref_3109_load_0_ack_1 : boolean;
  signal type_cast_3522_inst_req_1 : boolean;
  signal type_cast_3123_inst_req_0 : boolean;
  signal if_stmt_3486_branch_ack_0 : boolean;
  signal type_cast_3123_inst_ack_0 : boolean;
  signal type_cast_3123_inst_req_1 : boolean;
  signal type_cast_3123_inst_ack_1 : boolean;
  signal if_stmt_3512_branch_req_0 : boolean;
  signal type_cast_3498_inst_ack_1 : boolean;
  signal array_obj_ref_3567_index_offset_req_0 : boolean;
  signal array_obj_ref_3129_index_offset_req_0 : boolean;
  signal array_obj_ref_3129_index_offset_ack_0 : boolean;
  signal type_cast_3348_inst_req_0 : boolean;
  signal array_obj_ref_3129_index_offset_req_1 : boolean;
  signal if_stmt_3486_branch_ack_1 : boolean;
  signal array_obj_ref_3129_index_offset_ack_1 : boolean;
  signal addr_of_3130_final_reg_req_0 : boolean;
  signal addr_of_3130_final_reg_ack_0 : boolean;
  signal if_stmt_3486_branch_req_0 : boolean;
  signal addr_of_3130_final_reg_req_1 : boolean;
  signal addr_of_3130_final_reg_ack_1 : boolean;
  signal type_cast_3498_inst_req_1 : boolean;
  signal type_cast_3498_inst_ack_0 : boolean;
  signal type_cast_3498_inst_req_0 : boolean;
  signal type_cast_3335_inst_ack_1 : boolean;
  signal type_cast_3352_inst_req_0 : boolean;
  signal ptr_deref_3133_store_0_req_0 : boolean;
  signal if_stmt_3429_branch_ack_0 : boolean;
  signal ptr_deref_3133_store_0_ack_0 : boolean;
  signal type_cast_3441_inst_ack_1 : boolean;
  signal type_cast_3335_inst_req_1 : boolean;
  signal ptr_deref_3133_store_0_req_1 : boolean;
  signal ptr_deref_3133_store_0_ack_1 : boolean;
  signal addr_of_3568_final_reg_ack_1 : boolean;
  signal addr_of_4177_final_reg_req_1 : boolean;
  signal addr_of_3568_final_reg_req_1 : boolean;
  signal type_cast_3522_inst_ack_0 : boolean;
  signal type_cast_3141_inst_req_0 : boolean;
  signal type_cast_3141_inst_ack_0 : boolean;
  signal type_cast_3441_inst_req_1 : boolean;
  signal type_cast_3561_inst_ack_1 : boolean;
  signal type_cast_3141_inst_req_1 : boolean;
  signal type_cast_3141_inst_ack_1 : boolean;
  signal if_stmt_3429_branch_ack_1 : boolean;
  signal type_cast_3561_inst_req_1 : boolean;
  signal if_stmt_3156_branch_req_0 : boolean;
  signal type_cast_3335_inst_ack_0 : boolean;
  signal if_stmt_3156_branch_ack_1 : boolean;
  signal type_cast_3441_inst_ack_0 : boolean;
  signal type_cast_3335_inst_req_0 : boolean;
  signal if_stmt_3156_branch_ack_0 : boolean;
  signal type_cast_3441_inst_req_0 : boolean;
  signal addr_of_3568_final_reg_ack_0 : boolean;
  signal type_cast_3522_inst_req_0 : boolean;
  signal type_cast_3180_inst_req_0 : boolean;
  signal type_cast_3477_inst_ack_1 : boolean;
  signal type_cast_3180_inst_ack_0 : boolean;
  signal type_cast_3561_inst_ack_0 : boolean;
  signal type_cast_3561_inst_req_0 : boolean;
  signal type_cast_3180_inst_req_1 : boolean;
  signal type_cast_3477_inst_req_1 : boolean;
  signal type_cast_3180_inst_ack_1 : boolean;
  signal addr_of_3568_final_reg_req_0 : boolean;
  signal if_stmt_3429_branch_req_0 : boolean;
  signal LOAD_col_high_3183_load_0_req_0 : boolean;
  signal LOAD_col_high_3183_load_0_ack_0 : boolean;
  signal LOAD_col_high_3183_load_0_req_1 : boolean;
  signal LOAD_col_high_3183_load_0_ack_1 : boolean;
  signal type_cast_3420_inst_ack_1 : boolean;
  signal type_cast_3420_inst_req_1 : boolean;
  signal type_cast_3331_inst_ack_1 : boolean;
  signal type_cast_3187_inst_req_0 : boolean;
  signal type_cast_3187_inst_ack_0 : boolean;
  signal type_cast_3187_inst_req_1 : boolean;
  signal type_cast_3477_inst_ack_0 : boolean;
  signal type_cast_3187_inst_ack_1 : boolean;
  signal LOAD_col_high_3494_load_0_ack_1 : boolean;
  signal LOAD_col_high_3494_load_0_req_1 : boolean;
  signal type_cast_3477_inst_req_0 : boolean;
  signal type_cast_3207_inst_req_0 : boolean;
  signal type_cast_3207_inst_ack_0 : boolean;
  signal type_cast_3207_inst_req_1 : boolean;
  signal type_cast_3207_inst_ack_1 : boolean;
  signal type_cast_3527_inst_ack_1 : boolean;
  signal type_cast_3331_inst_req_1 : boolean;
  signal type_cast_3527_inst_req_1 : boolean;
  signal type_cast_3224_inst_req_0 : boolean;
  signal type_cast_3224_inst_ack_0 : boolean;
  signal type_cast_3224_inst_req_1 : boolean;
  signal type_cast_3224_inst_ack_1 : boolean;
  signal type_cast_3420_inst_ack_0 : boolean;
  signal type_cast_3420_inst_req_0 : boolean;
  signal type_cast_3348_inst_ack_1 : boolean;
  signal LOAD_row_high_3227_load_0_req_0 : boolean;
  signal LOAD_row_high_3227_load_0_ack_0 : boolean;
  signal type_cast_3348_inst_req_1 : boolean;
  signal LOAD_row_high_3227_load_0_req_1 : boolean;
  signal LOAD_row_high_3227_load_0_ack_1 : boolean;
  signal ptr_deref_3571_store_0_req_0 : boolean;
  signal type_cast_3527_inst_ack_0 : boolean;
  signal type_cast_3527_inst_req_0 : boolean;
  signal type_cast_3231_inst_req_0 : boolean;
  signal type_cast_3231_inst_ack_0 : boolean;
  signal type_cast_3231_inst_req_1 : boolean;
  signal type_cast_3231_inst_ack_1 : boolean;
  signal array_obj_ref_3567_index_offset_ack_1 : boolean;
  signal if_stmt_3255_branch_req_0 : boolean;
  signal if_stmt_3255_branch_ack_1 : boolean;
  signal if_stmt_3255_branch_ack_0 : boolean;
  signal LOAD_row_high_3437_load_0_ack_1 : boolean;
  signal if_stmt_3467_branch_ack_0 : boolean;
  signal type_cast_3299_inst_req_0 : boolean;
  signal type_cast_3299_inst_ack_0 : boolean;
  signal LOAD_row_high_3437_load_0_req_1 : boolean;
  signal type_cast_3299_inst_req_1 : boolean;
  signal type_cast_3299_inst_ack_1 : boolean;
  signal LOAD_col_high_3494_load_0_ack_0 : boolean;
  signal type_cast_3309_inst_req_0 : boolean;
  signal type_cast_3309_inst_ack_0 : boolean;
  signal type_cast_3973_inst_ack_1 : boolean;
  signal type_cast_3309_inst_req_1 : boolean;
  signal type_cast_3309_inst_ack_1 : boolean;
  signal type_cast_3883_inst_ack_1 : boolean;
  signal LOAD_pad_3318_load_0_req_0 : boolean;
  signal LOAD_pad_3318_load_0_ack_0 : boolean;
  signal LOAD_pad_3318_load_0_req_1 : boolean;
  signal LOAD_pad_3318_load_0_ack_1 : boolean;
  signal type_cast_4018_inst_req_0 : boolean;
  signal LOAD_row_high_3969_load_0_req_0 : boolean;
  signal LOAD_row_high_3969_load_0_ack_0 : boolean;
  signal type_cast_4048_inst_req_1 : boolean;
  signal type_cast_4170_inst_ack_1 : boolean;
  signal LOAD_depth_high_3321_load_0_req_0 : boolean;
  signal LOAD_depth_high_3321_load_0_ack_0 : boolean;
  signal type_cast_4018_inst_ack_0 : boolean;
  signal LOAD_depth_high_3321_load_0_req_1 : boolean;
  signal LOAD_depth_high_3321_load_0_ack_1 : boolean;
  signal type_cast_4018_inst_req_1 : boolean;
  signal type_cast_4018_inst_ack_1 : boolean;
  signal LOAD_out_depth_high_3324_load_0_req_0 : boolean;
  signal LOAD_out_depth_high_3324_load_0_ack_0 : boolean;
  signal LOAD_out_depth_high_3324_load_0_req_1 : boolean;
  signal LOAD_out_depth_high_3324_load_0_ack_1 : boolean;
  signal LOAD_out_col_high_3327_load_0_req_0 : boolean;
  signal LOAD_out_col_high_3327_load_0_ack_0 : boolean;
  signal LOAD_out_col_high_3327_load_0_req_1 : boolean;
  signal LOAD_out_col_high_3327_load_0_ack_1 : boolean;
  signal type_cast_3331_inst_req_0 : boolean;
  signal type_cast_3331_inst_ack_0 : boolean;
  signal ptr_deref_3571_store_0_ack_0 : boolean;
  signal ptr_deref_3571_store_0_req_1 : boolean;
  signal ptr_deref_3571_store_0_ack_1 : boolean;
  signal type_cast_3580_inst_req_0 : boolean;
  signal type_cast_3580_inst_ack_0 : boolean;
  signal type_cast_3580_inst_req_1 : boolean;
  signal type_cast_3580_inst_ack_1 : boolean;
  signal type_cast_3644_inst_req_0 : boolean;
  signal type_cast_3644_inst_ack_0 : boolean;
  signal type_cast_3644_inst_req_1 : boolean;
  signal type_cast_3644_inst_ack_1 : boolean;
  signal array_obj_ref_3650_index_offset_req_0 : boolean;
  signal array_obj_ref_3650_index_offset_ack_0 : boolean;
  signal array_obj_ref_3650_index_offset_req_1 : boolean;
  signal array_obj_ref_3650_index_offset_ack_1 : boolean;
  signal addr_of_3651_final_reg_req_0 : boolean;
  signal addr_of_3651_final_reg_ack_0 : boolean;
  signal addr_of_3651_final_reg_req_1 : boolean;
  signal addr_of_3651_final_reg_ack_1 : boolean;
  signal array_obj_ref_4176_index_offset_req_1 : boolean;
  signal type_cast_4048_inst_req_0 : boolean;
  signal type_cast_3973_inst_req_1 : boolean;
  signal ptr_deref_3655_load_0_req_0 : boolean;
  signal ptr_deref_3655_load_0_ack_0 : boolean;
  signal if_stmt_3961_branch_ack_0 : boolean;
  signal type_cast_3973_inst_ack_0 : boolean;
  signal ptr_deref_3655_load_0_req_1 : boolean;
  signal ptr_deref_3655_load_0_ack_1 : boolean;
  signal array_obj_ref_4176_index_offset_ack_0 : boolean;
  signal addr_of_4094_final_reg_ack_1 : boolean;
  signal LOAD_col_high_4014_load_0_ack_1 : boolean;
  signal type_cast_3883_inst_req_1 : boolean;
  signal LOAD_col_high_4014_load_0_req_1 : boolean;
  signal type_cast_3669_inst_req_0 : boolean;
  signal type_cast_3669_inst_ack_0 : boolean;
  signal type_cast_3669_inst_req_1 : boolean;
  signal type_cast_3669_inst_ack_1 : boolean;
  signal array_obj_ref_4176_index_offset_req_0 : boolean;
  signal addr_of_4705_final_reg_ack_1 : boolean;
  signal addr_of_4094_final_reg_req_1 : boolean;
  signal addr_of_4094_final_reg_ack_0 : boolean;
  signal addr_of_4094_final_reg_req_0 : boolean;
  signal type_cast_4170_inst_req_1 : boolean;
  signal array_obj_ref_3675_index_offset_req_0 : boolean;
  signal array_obj_ref_3675_index_offset_ack_0 : boolean;
  signal array_obj_ref_3675_index_offset_req_1 : boolean;
  signal array_obj_ref_3675_index_offset_ack_1 : boolean;
  signal type_cast_4087_inst_ack_1 : boolean;
  signal if_stmt_3961_branch_ack_1 : boolean;
  signal type_cast_4087_inst_req_1 : boolean;
  signal addr_of_3676_final_reg_req_0 : boolean;
  signal addr_of_3676_final_reg_ack_0 : boolean;
  signal addr_of_3676_final_reg_req_1 : boolean;
  signal addr_of_3676_final_reg_ack_1 : boolean;
  signal if_stmt_3961_branch_req_0 : boolean;
  signal array_obj_ref_4093_index_offset_ack_1 : boolean;
  signal array_obj_ref_4093_index_offset_req_1 : boolean;
  signal LOAD_col_high_4014_load_0_ack_0 : boolean;
  signal type_cast_4087_inst_ack_0 : boolean;
  signal LOAD_col_high_4014_load_0_req_0 : boolean;
  signal type_cast_3973_inst_req_0 : boolean;
  signal type_cast_4087_inst_req_0 : boolean;
  signal ptr_deref_3679_store_0_req_0 : boolean;
  signal ptr_deref_3679_store_0_ack_0 : boolean;
  signal ptr_deref_3679_store_0_req_1 : boolean;
  signal ptr_deref_3679_store_0_ack_1 : boolean;
  signal type_cast_4170_inst_ack_0 : boolean;
  signal ptr_deref_4097_store_0_ack_1 : boolean;
  signal type_cast_3687_inst_req_0 : boolean;
  signal type_cast_3687_inst_ack_0 : boolean;
  signal ptr_deref_4097_store_0_req_1 : boolean;
  signal type_cast_3687_inst_req_1 : boolean;
  signal type_cast_3687_inst_ack_1 : boolean;
  signal if_stmt_3702_branch_req_0 : boolean;
  signal type_cast_4170_inst_req_0 : boolean;
  signal type_cast_3952_inst_ack_1 : boolean;
  signal if_stmt_3702_branch_ack_1 : boolean;
  signal type_cast_3952_inst_req_1 : boolean;
  signal if_stmt_3702_branch_ack_0 : boolean;
  signal if_stmt_4038_branch_ack_0 : boolean;
  signal array_obj_ref_4093_index_offset_ack_0 : boolean;
  signal type_cast_3726_inst_req_0 : boolean;
  signal type_cast_3726_inst_ack_0 : boolean;
  signal type_cast_3726_inst_req_1 : boolean;
  signal type_cast_3726_inst_ack_1 : boolean;
  signal LOAD_col_high_3729_load_0_req_0 : boolean;
  signal LOAD_col_high_3729_load_0_ack_0 : boolean;
  signal LOAD_col_high_3729_load_0_req_1 : boolean;
  signal LOAD_col_high_3729_load_0_ack_1 : boolean;
  signal array_obj_ref_4093_index_offset_req_0 : boolean;
  signal type_cast_3883_inst_ack_0 : boolean;
  signal ptr_deref_4097_store_0_ack_0 : boolean;
  signal type_cast_3733_inst_req_0 : boolean;
  signal type_cast_4053_inst_ack_1 : boolean;
  signal type_cast_3733_inst_ack_0 : boolean;
  signal if_stmt_4038_branch_ack_1 : boolean;
  signal ptr_deref_4097_store_0_req_0 : boolean;
  signal type_cast_3733_inst_req_1 : boolean;
  signal type_cast_4053_inst_req_1 : boolean;
  signal type_cast_3733_inst_ack_1 : boolean;
  signal type_cast_3747_inst_req_0 : boolean;
  signal type_cast_3747_inst_ack_0 : boolean;
  signal type_cast_3747_inst_req_1 : boolean;
  signal type_cast_4053_inst_ack_0 : boolean;
  signal type_cast_3747_inst_ack_1 : boolean;
  signal type_cast_3883_inst_req_0 : boolean;
  signal type_cast_4053_inst_req_0 : boolean;
  signal type_cast_3763_inst_req_0 : boolean;
  signal type_cast_3763_inst_ack_0 : boolean;
  signal type_cast_3763_inst_req_1 : boolean;
  signal type_cast_3763_inst_ack_1 : boolean;
  signal if_stmt_4006_branch_ack_0 : boolean;
  signal if_stmt_4006_branch_ack_1 : boolean;
  signal LOAD_row_high_3766_load_0_req_0 : boolean;
  signal LOAD_row_high_3766_load_0_ack_0 : boolean;
  signal LOAD_row_high_3766_load_0_req_1 : boolean;
  signal LOAD_row_high_3766_load_0_ack_1 : boolean;
  signal if_stmt_4006_branch_req_0 : boolean;
  signal addr_of_4177_final_reg_ack_0 : boolean;
  signal type_cast_3770_inst_req_0 : boolean;
  signal type_cast_3770_inst_ack_0 : boolean;
  signal if_stmt_4038_branch_req_0 : boolean;
  signal type_cast_3770_inst_req_1 : boolean;
  signal type_cast_3770_inst_ack_1 : boolean;
  signal type_cast_3952_inst_ack_0 : boolean;
  signal type_cast_3952_inst_req_0 : boolean;
  signal addr_of_4177_final_reg_req_0 : boolean;
  signal if_stmt_3794_branch_req_0 : boolean;
  signal if_stmt_3794_branch_ack_1 : boolean;
  signal if_stmt_3794_branch_ack_0 : boolean;
  signal type_cast_3834_inst_req_0 : boolean;
  signal type_cast_3834_inst_ack_0 : boolean;
  signal type_cast_3834_inst_req_1 : boolean;
  signal type_cast_3834_inst_ack_1 : boolean;
  signal array_obj_ref_4176_index_offset_ack_1 : boolean;
  signal type_cast_4048_inst_ack_1 : boolean;
  signal LOAD_pad_3849_load_0_req_0 : boolean;
  signal LOAD_pad_3849_load_0_ack_0 : boolean;
  signal LOAD_row_high_3969_load_0_ack_1 : boolean;
  signal LOAD_pad_3849_load_0_req_1 : boolean;
  signal type_cast_3997_inst_ack_1 : boolean;
  signal LOAD_pad_3849_load_0_ack_1 : boolean;
  signal type_cast_3997_inst_req_1 : boolean;
  signal addr_of_4705_final_reg_req_1 : boolean;
  signal type_cast_3997_inst_ack_0 : boolean;
  signal type_cast_3997_inst_req_0 : boolean;
  signal LOAD_row_high_3969_load_0_req_1 : boolean;
  signal LOAD_depth_high_3852_load_0_req_0 : boolean;
  signal LOAD_depth_high_3852_load_0_ack_0 : boolean;
  signal LOAD_depth_high_3852_load_0_req_1 : boolean;
  signal LOAD_depth_high_3852_load_0_ack_1 : boolean;
  signal type_cast_4106_inst_ack_1 : boolean;
  signal type_cast_4106_inst_req_1 : boolean;
  signal if_stmt_3987_branch_ack_0 : boolean;
  signal LOAD_out_depth_high_3855_load_0_req_0 : boolean;
  signal LOAD_out_depth_high_3855_load_0_ack_0 : boolean;
  signal if_stmt_3987_branch_ack_1 : boolean;
  signal LOAD_out_depth_high_3855_load_0_req_1 : boolean;
  signal LOAD_out_depth_high_3855_load_0_ack_1 : boolean;
  signal type_cast_4106_inst_ack_0 : boolean;
  signal if_stmt_3987_branch_req_0 : boolean;
  signal addr_of_4177_final_reg_ack_1 : boolean;
  signal LOAD_out_col_high_3858_load_0_req_0 : boolean;
  signal LOAD_out_col_high_3858_load_0_ack_0 : boolean;
  signal LOAD_out_col_high_3858_load_0_req_1 : boolean;
  signal LOAD_out_col_high_3858_load_0_ack_1 : boolean;
  signal type_cast_4106_inst_req_0 : boolean;
  signal type_cast_3862_inst_req_0 : boolean;
  signal ptr_deref_4625_store_0_req_0 : boolean;
  signal type_cast_3862_inst_ack_0 : boolean;
  signal type_cast_3862_inst_req_1 : boolean;
  signal type_cast_3862_inst_ack_1 : boolean;
  signal ptr_deref_4625_store_0_ack_0 : boolean;
  signal type_cast_3866_inst_req_0 : boolean;
  signal type_cast_3866_inst_ack_0 : boolean;
  signal ptr_deref_4709_load_0_req_1 : boolean;
  signal type_cast_3866_inst_req_1 : boolean;
  signal type_cast_3866_inst_ack_1 : boolean;
  signal type_cast_3870_inst_req_0 : boolean;
  signal type_cast_3870_inst_ack_0 : boolean;
  signal type_cast_3870_inst_req_1 : boolean;
  signal type_cast_3870_inst_ack_1 : boolean;
  signal type_cast_3879_inst_req_0 : boolean;
  signal type_cast_3879_inst_ack_0 : boolean;
  signal type_cast_3879_inst_req_1 : boolean;
  signal type_cast_3879_inst_ack_1 : boolean;
  signal ptr_deref_4181_load_0_req_0 : boolean;
  signal ptr_deref_4181_load_0_ack_0 : boolean;
  signal ptr_deref_4181_load_0_req_1 : boolean;
  signal ptr_deref_4181_load_0_ack_1 : boolean;
  signal type_cast_4195_inst_req_0 : boolean;
  signal type_cast_4195_inst_ack_0 : boolean;
  signal type_cast_4195_inst_req_1 : boolean;
  signal type_cast_4195_inst_ack_1 : boolean;
  signal addr_of_4705_final_reg_ack_0 : boolean;
  signal addr_of_4705_final_reg_req_0 : boolean;
  signal type_cast_4581_inst_ack_1 : boolean;
  signal type_cast_4581_inst_req_1 : boolean;
  signal array_obj_ref_4201_index_offset_req_0 : boolean;
  signal array_obj_ref_4201_index_offset_ack_0 : boolean;
  signal array_obj_ref_4201_index_offset_req_1 : boolean;
  signal array_obj_ref_4201_index_offset_ack_1 : boolean;
  signal type_cast_4581_inst_ack_0 : boolean;
  signal type_cast_4581_inst_req_0 : boolean;
  signal addr_of_4202_final_reg_req_0 : boolean;
  signal addr_of_4202_final_reg_ack_0 : boolean;
  signal addr_of_4202_final_reg_req_1 : boolean;
  signal addr_of_4202_final_reg_ack_1 : boolean;
  signal type_cast_4576_inst_ack_1 : boolean;
  signal ptr_deref_4205_store_0_req_0 : boolean;
  signal ptr_deref_4205_store_0_ack_0 : boolean;
  signal type_cast_4576_inst_req_1 : boolean;
  signal ptr_deref_4205_store_0_req_1 : boolean;
  signal ptr_deref_4205_store_0_ack_1 : boolean;
  signal type_cast_4723_inst_ack_0 : boolean;
  signal type_cast_4723_inst_req_0 : boolean;
  signal ptr_deref_4709_load_0_ack_0 : boolean;
  signal type_cast_4213_inst_req_0 : boolean;
  signal type_cast_4213_inst_ack_0 : boolean;
  signal ptr_deref_4709_load_0_req_0 : boolean;
  signal type_cast_4213_inst_req_1 : boolean;
  signal type_cast_4213_inst_ack_1 : boolean;
  signal if_stmt_4228_branch_req_0 : boolean;
  signal type_cast_4576_inst_ack_0 : boolean;
  signal if_stmt_4228_branch_ack_1 : boolean;
  signal ptr_deref_4625_store_0_ack_1 : boolean;
  signal type_cast_4576_inst_req_0 : boolean;
  signal if_stmt_4228_branch_ack_0 : boolean;
  signal ptr_deref_4625_store_0_req_1 : boolean;
  signal array_obj_ref_4704_index_offset_ack_1 : boolean;
  signal type_cast_4698_inst_ack_1 : boolean;
  signal type_cast_4698_inst_req_1 : boolean;
  signal type_cast_4252_inst_req_0 : boolean;
  signal type_cast_4252_inst_ack_0 : boolean;
  signal type_cast_4252_inst_req_1 : boolean;
  signal type_cast_4252_inst_ack_1 : boolean;
  signal array_obj_ref_4704_index_offset_req_1 : boolean;
  signal LOAD_col_high_4255_load_0_req_0 : boolean;
  signal LOAD_col_high_4255_load_0_ack_0 : boolean;
  signal LOAD_col_high_4255_load_0_req_1 : boolean;
  signal LOAD_col_high_4255_load_0_ack_1 : boolean;
  signal type_cast_4259_inst_req_0 : boolean;
  signal type_cast_4698_inst_ack_0 : boolean;
  signal type_cast_4259_inst_ack_0 : boolean;
  signal if_stmt_4566_branch_ack_0 : boolean;
  signal type_cast_4259_inst_req_1 : boolean;
  signal type_cast_4698_inst_req_0 : boolean;
  signal type_cast_4259_inst_ack_1 : boolean;
  signal array_obj_ref_4704_index_offset_ack_0 : boolean;
  signal type_cast_4279_inst_req_0 : boolean;
  signal type_cast_4279_inst_ack_0 : boolean;
  signal type_cast_4279_inst_req_1 : boolean;
  signal type_cast_4279_inst_ack_1 : boolean;
  signal array_obj_ref_4704_index_offset_req_0 : boolean;
  signal addr_of_4622_final_reg_ack_1 : boolean;
  signal addr_of_4622_final_reg_req_1 : boolean;
  signal type_cast_4296_inst_req_0 : boolean;
  signal type_cast_4296_inst_ack_0 : boolean;
  signal type_cast_4296_inst_req_1 : boolean;
  signal type_cast_4296_inst_ack_1 : boolean;
  signal type_cast_1674_inst_ack_1 : boolean;
  signal type_cast_4615_inst_ack_1 : boolean;
  signal type_cast_4615_inst_req_1 : boolean;
  signal addr_of_4622_final_reg_ack_0 : boolean;
  signal addr_of_4622_final_reg_req_0 : boolean;
  signal LOAD_row_high_4299_load_0_req_0 : boolean;
  signal LOAD_row_high_4299_load_0_ack_0 : boolean;
  signal LOAD_row_high_4299_load_0_req_1 : boolean;
  signal LOAD_row_high_4299_load_0_ack_1 : boolean;
  signal ptr_deref_4709_load_0_ack_1 : boolean;
  signal if_stmt_4566_branch_ack_1 : boolean;
  signal array_obj_ref_4621_index_offset_ack_1 : boolean;
  signal array_obj_ref_4621_index_offset_req_1 : boolean;
  signal type_cast_4634_inst_ack_1 : boolean;
  signal type_cast_4303_inst_req_0 : boolean;
  signal type_cast_4634_inst_req_1 : boolean;
  signal type_cast_4303_inst_ack_0 : boolean;
  signal type_cast_4303_inst_req_1 : boolean;
  signal type_cast_4303_inst_ack_1 : boolean;
  signal type_cast_4615_inst_ack_0 : boolean;
  signal if_stmt_4315_branch_req_0 : boolean;
  signal if_stmt_4315_branch_ack_1 : boolean;
  signal if_stmt_4315_branch_ack_0 : boolean;
  signal array_obj_ref_4621_index_offset_ack_0 : boolean;
  signal type_cast_4359_inst_req_0 : boolean;
  signal type_cast_4634_inst_ack_0 : boolean;
  signal type_cast_4359_inst_ack_0 : boolean;
  signal type_cast_4359_inst_req_1 : boolean;
  signal type_cast_4634_inst_req_0 : boolean;
  signal type_cast_4359_inst_ack_1 : boolean;
  signal type_cast_4615_inst_req_0 : boolean;
  signal array_obj_ref_4621_index_offset_req_0 : boolean;
  signal type_cast_4369_inst_req_0 : boolean;
  signal type_cast_4369_inst_ack_0 : boolean;
  signal type_cast_4369_inst_req_1 : boolean;
  signal type_cast_4369_inst_ack_1 : boolean;
  signal type_cast_1800_inst_ack_1 : boolean;
  signal phi_stmt_1669_req_1 : boolean;
  signal LOAD_pad_4384_load_0_req_0 : boolean;
  signal LOAD_pad_4384_load_0_ack_0 : boolean;
  signal LOAD_pad_4384_load_0_req_1 : boolean;
  signal LOAD_pad_4384_load_0_ack_1 : boolean;
  signal phi_stmt_1675_ack_0 : boolean;
  signal type_cast_1694_inst_ack_1 : boolean;
  signal LOAD_depth_high_4387_load_0_req_0 : boolean;
  signal LOAD_depth_high_4387_load_0_ack_0 : boolean;
  signal LOAD_depth_high_4387_load_0_req_1 : boolean;
  signal LOAD_depth_high_4387_load_0_ack_1 : boolean;
  signal type_cast_1680_inst_req_0 : boolean;
  signal LOAD_out_depth_high_4390_load_0_req_0 : boolean;
  signal LOAD_out_depth_high_4390_load_0_ack_0 : boolean;
  signal LOAD_out_depth_high_4390_load_0_req_1 : boolean;
  signal LOAD_out_depth_high_4390_load_0_ack_1 : boolean;
  signal phi_stmt_1681_ack_0 : boolean;
  signal LOAD_out_col_high_4393_load_0_req_0 : boolean;
  signal LOAD_out_col_high_4393_load_0_ack_0 : boolean;
  signal type_cast_1680_inst_ack_0 : boolean;
  signal LOAD_out_col_high_4393_load_0_req_1 : boolean;
  signal LOAD_out_col_high_4393_load_0_ack_1 : boolean;
  signal type_cast_4397_inst_req_0 : boolean;
  signal type_cast_4397_inst_ack_0 : boolean;
  signal type_cast_4397_inst_req_1 : boolean;
  signal type_cast_4397_inst_ack_1 : boolean;
  signal type_cast_1809_inst_req_0 : boolean;
  signal type_cast_4401_inst_req_0 : boolean;
  signal type_cast_4401_inst_ack_0 : boolean;
  signal type_cast_1793_inst_req_1 : boolean;
  signal type_cast_4401_inst_req_1 : boolean;
  signal type_cast_4401_inst_ack_1 : boolean;
  signal type_cast_1680_inst_req_1 : boolean;
  signal type_cast_1793_inst_ack_1 : boolean;
  signal type_cast_4405_inst_req_0 : boolean;
  signal type_cast_4405_inst_ack_0 : boolean;
  signal type_cast_4405_inst_req_1 : boolean;
  signal type_cast_1680_inst_ack_1 : boolean;
  signal type_cast_4405_inst_ack_1 : boolean;
  signal type_cast_1809_inst_ack_0 : boolean;
  signal phi_stmt_1790_req_0 : boolean;
  signal type_cast_4414_inst_req_0 : boolean;
  signal phi_stmt_1691_req_0 : boolean;
  signal type_cast_4414_inst_ack_0 : boolean;
  signal type_cast_4414_inst_req_1 : boolean;
  signal type_cast_4414_inst_ack_1 : boolean;
  signal phi_stmt_1675_req_1 : boolean;
  signal type_cast_4418_inst_req_0 : boolean;
  signal type_cast_4418_inst_ack_0 : boolean;
  signal type_cast_4418_inst_req_1 : boolean;
  signal type_cast_4418_inst_ack_1 : boolean;
  signal type_cast_4486_inst_req_0 : boolean;
  signal type_cast_4486_inst_ack_0 : boolean;
  signal type_cast_4486_inst_req_1 : boolean;
  signal type_cast_4486_inst_ack_1 : boolean;
  signal phi_stmt_1797_req_0 : boolean;
  signal if_stmt_4495_branch_req_0 : boolean;
  signal if_stmt_4495_branch_ack_1 : boolean;
  signal if_stmt_4495_branch_ack_0 : boolean;
  signal LOAD_row_high_4503_load_0_req_0 : boolean;
  signal LOAD_row_high_4503_load_0_ack_0 : boolean;
  signal LOAD_row_high_4503_load_0_req_1 : boolean;
  signal LOAD_row_high_4503_load_0_ack_1 : boolean;
  signal type_cast_4507_inst_req_0 : boolean;
  signal type_cast_4507_inst_ack_0 : boolean;
  signal type_cast_4507_inst_req_1 : boolean;
  signal type_cast_4507_inst_ack_1 : boolean;
  signal if_stmt_4521_branch_req_0 : boolean;
  signal if_stmt_4521_branch_ack_1 : boolean;
  signal if_stmt_4521_branch_ack_0 : boolean;
  signal type_cast_4531_inst_req_0 : boolean;
  signal type_cast_4531_inst_ack_0 : boolean;
  signal type_cast_4531_inst_req_1 : boolean;
  signal type_cast_4531_inst_ack_1 : boolean;
  signal if_stmt_4540_branch_req_0 : boolean;
  signal if_stmt_4540_branch_ack_1 : boolean;
  signal if_stmt_4540_branch_ack_0 : boolean;
  signal LOAD_col_high_4548_load_0_req_0 : boolean;
  signal LOAD_col_high_4548_load_0_ack_0 : boolean;
  signal LOAD_col_high_4548_load_0_req_1 : boolean;
  signal LOAD_col_high_4548_load_0_ack_1 : boolean;
  signal type_cast_4552_inst_req_0 : boolean;
  signal type_cast_4552_inst_ack_0 : boolean;
  signal type_cast_4552_inst_req_1 : boolean;
  signal type_cast_4552_inst_ack_1 : boolean;
  signal if_stmt_4566_branch_req_0 : boolean;
  signal type_cast_4723_inst_req_1 : boolean;
  signal type_cast_4723_inst_ack_1 : boolean;
  signal array_obj_ref_4729_index_offset_req_0 : boolean;
  signal array_obj_ref_4729_index_offset_ack_0 : boolean;
  signal array_obj_ref_4729_index_offset_req_1 : boolean;
  signal array_obj_ref_4729_index_offset_ack_1 : boolean;
  signal addr_of_4730_final_reg_req_0 : boolean;
  signal addr_of_4730_final_reg_ack_0 : boolean;
  signal addr_of_4730_final_reg_req_1 : boolean;
  signal addr_of_4730_final_reg_ack_1 : boolean;
  signal ptr_deref_4733_store_0_req_0 : boolean;
  signal ptr_deref_4733_store_0_ack_0 : boolean;
  signal ptr_deref_4733_store_0_req_1 : boolean;
  signal ptr_deref_4733_store_0_ack_1 : boolean;
  signal type_cast_4741_inst_req_0 : boolean;
  signal type_cast_4741_inst_ack_0 : boolean;
  signal type_cast_4741_inst_req_1 : boolean;
  signal type_cast_4741_inst_ack_1 : boolean;
  signal if_stmt_4756_branch_req_0 : boolean;
  signal if_stmt_4756_branch_ack_1 : boolean;
  signal if_stmt_4756_branch_ack_0 : boolean;
  signal type_cast_4780_inst_req_0 : boolean;
  signal type_cast_4780_inst_ack_0 : boolean;
  signal type_cast_4780_inst_req_1 : boolean;
  signal type_cast_4780_inst_ack_1 : boolean;
  signal LOAD_col_high_4783_load_0_req_0 : boolean;
  signal LOAD_col_high_4783_load_0_ack_0 : boolean;
  signal LOAD_col_high_4783_load_0_req_1 : boolean;
  signal LOAD_col_high_4783_load_0_ack_1 : boolean;
  signal type_cast_1694_inst_req_1 : boolean;
  signal type_cast_1793_inst_ack_0 : boolean;
  signal type_cast_4787_inst_req_0 : boolean;
  signal type_cast_4787_inst_ack_0 : boolean;
  signal phi_stmt_1669_ack_0 : boolean;
  signal type_cast_1793_inst_req_0 : boolean;
  signal type_cast_4787_inst_req_1 : boolean;
  signal type_cast_1694_inst_ack_0 : boolean;
  signal type_cast_4787_inst_ack_1 : boolean;
  signal type_cast_1800_inst_req_1 : boolean;
  signal type_cast_1694_inst_req_0 : boolean;
  signal type_cast_4801_inst_req_0 : boolean;
  signal type_cast_4801_inst_ack_0 : boolean;
  signal type_cast_4801_inst_req_1 : boolean;
  signal type_cast_4801_inst_ack_1 : boolean;
  signal type_cast_1800_inst_ack_0 : boolean;
  signal type_cast_4817_inst_req_0 : boolean;
  signal type_cast_4817_inst_ack_0 : boolean;
  signal type_cast_4817_inst_req_1 : boolean;
  signal type_cast_4817_inst_ack_1 : boolean;
  signal phi_stmt_1681_req_1 : boolean;
  signal LOAD_row_high_4820_load_0_req_0 : boolean;
  signal LOAD_row_high_4820_load_0_ack_0 : boolean;
  signal LOAD_row_high_4820_load_0_req_1 : boolean;
  signal LOAD_row_high_4820_load_0_ack_1 : boolean;
  signal phi_stmt_1695_ack_0 : boolean;
  signal type_cast_4824_inst_req_0 : boolean;
  signal type_cast_4824_inst_ack_0 : boolean;
  signal phi_stmt_1669_req_0 : boolean;
  signal type_cast_4824_inst_req_1 : boolean;
  signal type_cast_4824_inst_ack_1 : boolean;
  signal type_cast_1800_inst_req_0 : boolean;
  signal type_cast_1672_inst_ack_1 : boolean;
  signal phi_stmt_1797_req_1 : boolean;
  signal if_stmt_4836_branch_req_0 : boolean;
  signal phi_stmt_1803_req_0 : boolean;
  signal type_cast_1672_inst_req_1 : boolean;
  signal if_stmt_4836_branch_ack_1 : boolean;
  signal if_stmt_4836_branch_ack_0 : boolean;
  signal type_cast_1809_inst_ack_1 : boolean;
  signal type_cast_1674_inst_req_1 : boolean;
  signal type_cast_1809_inst_req_1 : boolean;
  signal type_cast_1672_inst_ack_0 : boolean;
  signal phi_stmt_1691_ack_0 : boolean;
  signal type_cast_1802_inst_ack_1 : boolean;
  signal call_stmt_4866_call_req_0 : boolean;
  signal phi_stmt_1695_req_0 : boolean;
  signal call_stmt_4866_call_ack_0 : boolean;
  signal type_cast_1672_inst_req_0 : boolean;
  signal type_cast_1802_inst_req_1 : boolean;
  signal call_stmt_4866_call_req_1 : boolean;
  signal type_cast_1698_inst_ack_1 : boolean;
  signal call_stmt_4866_call_ack_1 : boolean;
  signal phi_stmt_747_req_0 : boolean;
  signal phi_stmt_1675_req_0 : boolean;
  signal phi_stmt_754_req_0 : boolean;
  signal phi_stmt_761_req_0 : boolean;
  signal type_cast_1698_inst_req_1 : boolean;
  signal type_cast_753_inst_req_0 : boolean;
  signal type_cast_753_inst_ack_0 : boolean;
  signal type_cast_753_inst_req_1 : boolean;
  signal type_cast_753_inst_ack_1 : boolean;
  signal phi_stmt_747_req_1 : boolean;
  signal type_cast_760_inst_req_0 : boolean;
  signal type_cast_760_inst_ack_0 : boolean;
  signal type_cast_1698_inst_ack_0 : boolean;
  signal type_cast_760_inst_req_1 : boolean;
  signal type_cast_760_inst_ack_1 : boolean;
  signal phi_stmt_754_req_1 : boolean;
  signal type_cast_1698_inst_req_0 : boolean;
  signal type_cast_767_inst_req_0 : boolean;
  signal type_cast_767_inst_ack_0 : boolean;
  signal type_cast_767_inst_req_1 : boolean;
  signal type_cast_767_inst_ack_1 : boolean;
  signal phi_stmt_761_req_1 : boolean;
  signal phi_stmt_1681_req_0 : boolean;
  signal phi_stmt_747_ack_0 : boolean;
  signal phi_stmt_754_ack_0 : boolean;
  signal phi_stmt_761_ack_0 : boolean;
  signal type_cast_1678_inst_ack_1 : boolean;
  signal type_cast_1684_inst_ack_1 : boolean;
  signal type_cast_1684_inst_req_1 : boolean;
  signal type_cast_1678_inst_req_1 : boolean;
  signal type_cast_1802_inst_ack_0 : boolean;
  signal type_cast_1678_inst_ack_0 : boolean;
  signal type_cast_1684_inst_ack_0 : boolean;
  signal type_cast_1684_inst_req_0 : boolean;
  signal type_cast_3813_inst_req_0 : boolean;
  signal type_cast_1802_inst_req_0 : boolean;
  signal type_cast_1678_inst_req_0 : boolean;
  signal type_cast_1674_inst_ack_0 : boolean;
  signal phi_stmt_1803_req_1 : boolean;
  signal type_cast_1674_inst_req_0 : boolean;
  signal type_cast_3813_inst_req_1 : boolean;
  signal type_cast_3813_inst_ack_1 : boolean;
  signal phi_stmt_3808_req_1 : boolean;
  signal type_cast_3804_inst_req_0 : boolean;
  signal type_cast_1160_inst_req_0 : boolean;
  signal type_cast_1160_inst_ack_0 : boolean;
  signal type_cast_1160_inst_req_1 : boolean;
  signal type_cast_1160_inst_ack_1 : boolean;
  signal type_cast_3409_inst_ack_0 : boolean;
  signal phi_stmt_1155_req_1 : boolean;
  signal type_cast_3804_inst_ack_0 : boolean;
  signal phi_stmt_3801_req_1 : boolean;
  signal type_cast_1166_inst_req_0 : boolean;
  signal type_cast_1166_inst_ack_0 : boolean;
  signal type_cast_1166_inst_req_1 : boolean;
  signal type_cast_1166_inst_ack_1 : boolean;
  signal phi_stmt_1161_req_1 : boolean;
  signal phi_stmt_1167_req_1 : boolean;
  signal type_cast_1158_inst_req_0 : boolean;
  signal type_cast_1158_inst_ack_0 : boolean;
  signal type_cast_1158_inst_req_1 : boolean;
  signal type_cast_1158_inst_ack_1 : boolean;
  signal phi_stmt_1155_req_0 : boolean;
  signal type_cast_1164_inst_req_0 : boolean;
  signal type_cast_1164_inst_ack_0 : boolean;
  signal type_cast_1164_inst_req_1 : boolean;
  signal type_cast_1164_inst_ack_1 : boolean;
  signal phi_stmt_1161_req_0 : boolean;
  signal type_cast_1170_inst_req_0 : boolean;
  signal type_cast_1170_inst_ack_0 : boolean;
  signal type_cast_1170_inst_req_1 : boolean;
  signal type_cast_1170_inst_ack_1 : boolean;
  signal phi_stmt_1167_req_0 : boolean;
  signal phi_stmt_1155_ack_0 : boolean;
  signal phi_stmt_1161_ack_0 : boolean;
  signal phi_stmt_1167_ack_0 : boolean;
  signal type_cast_1180_inst_req_0 : boolean;
  signal type_cast_1180_inst_ack_0 : boolean;
  signal type_cast_1180_inst_req_1 : boolean;
  signal type_cast_1180_inst_ack_1 : boolean;
  signal phi_stmt_1177_req_0 : boolean;
  signal type_cast_3409_inst_req_1 : boolean;
  signal type_cast_1184_inst_req_0 : boolean;
  signal type_cast_1184_inst_ack_0 : boolean;
  signal type_cast_3409_inst_ack_1 : boolean;
  signal type_cast_1184_inst_req_1 : boolean;
  signal type_cast_1184_inst_ack_1 : boolean;
  signal phi_stmt_1181_req_0 : boolean;
  signal phi_stmt_1177_ack_0 : boolean;
  signal phi_stmt_1181_ack_0 : boolean;
  signal type_cast_1281_inst_req_0 : boolean;
  signal type_cast_1281_inst_ack_0 : boolean;
  signal type_cast_1281_inst_req_1 : boolean;
  signal type_cast_1281_inst_ack_1 : boolean;
  signal phi_stmt_1276_req_1 : boolean;
  signal type_cast_1288_inst_req_0 : boolean;
  signal type_cast_1288_inst_ack_0 : boolean;
  signal type_cast_1288_inst_req_1 : boolean;
  signal type_cast_1288_inst_ack_1 : boolean;
  signal phi_stmt_1282_req_1 : boolean;
  signal type_cast_1295_inst_req_0 : boolean;
  signal type_cast_1295_inst_ack_0 : boolean;
  signal type_cast_1295_inst_req_1 : boolean;
  signal type_cast_1295_inst_ack_1 : boolean;
  signal phi_stmt_1289_req_1 : boolean;
  signal type_cast_1279_inst_req_0 : boolean;
  signal type_cast_1279_inst_ack_0 : boolean;
  signal type_cast_1279_inst_req_1 : boolean;
  signal type_cast_1279_inst_ack_1 : boolean;
  signal phi_stmt_1276_req_0 : boolean;
  signal phi_stmt_1282_req_0 : boolean;
  signal phi_stmt_1289_req_0 : boolean;
  signal phi_stmt_1276_ack_0 : boolean;
  signal phi_stmt_1282_ack_0 : boolean;
  signal phi_stmt_1289_ack_0 : boolean;
  signal phi_stmt_1790_req_1 : boolean;
  signal phi_stmt_1790_ack_0 : boolean;
  signal phi_stmt_1797_ack_0 : boolean;
  signal phi_stmt_1803_ack_0 : boolean;
  signal phi_stmt_2196_req_1 : boolean;
  signal type_cast_2206_inst_req_0 : boolean;
  signal type_cast_2206_inst_ack_0 : boolean;
  signal type_cast_2206_inst_req_1 : boolean;
  signal type_cast_2206_inst_ack_1 : boolean;
  signal phi_stmt_2203_req_0 : boolean;
  signal type_cast_2212_inst_req_0 : boolean;
  signal type_cast_2212_inst_ack_0 : boolean;
  signal type_cast_2212_inst_req_1 : boolean;
  signal type_cast_2212_inst_ack_1 : boolean;
  signal phi_stmt_2209_req_0 : boolean;
  signal type_cast_2199_inst_req_0 : boolean;
  signal type_cast_2199_inst_ack_0 : boolean;
  signal type_cast_2199_inst_req_1 : boolean;
  signal type_cast_2199_inst_ack_1 : boolean;
  signal phi_stmt_2196_req_0 : boolean;
  signal type_cast_2208_inst_req_0 : boolean;
  signal type_cast_2208_inst_ack_0 : boolean;
  signal type_cast_2208_inst_req_1 : boolean;
  signal type_cast_2208_inst_ack_1 : boolean;
  signal phi_stmt_2203_req_1 : boolean;
  signal type_cast_2214_inst_req_0 : boolean;
  signal type_cast_2214_inst_ack_0 : boolean;
  signal type_cast_2214_inst_req_1 : boolean;
  signal type_cast_2214_inst_ack_1 : boolean;
  signal phi_stmt_2209_req_1 : boolean;
  signal phi_stmt_2196_ack_0 : boolean;
  signal phi_stmt_2203_ack_0 : boolean;
  signal phi_stmt_2209_ack_0 : boolean;
  signal type_cast_2221_inst_req_0 : boolean;
  signal type_cast_2221_inst_ack_0 : boolean;
  signal type_cast_2221_inst_req_1 : boolean;
  signal type_cast_2221_inst_ack_1 : boolean;
  signal phi_stmt_2218_req_0 : boolean;
  signal type_cast_2225_inst_req_0 : boolean;
  signal type_cast_2225_inst_ack_0 : boolean;
  signal type_cast_2225_inst_req_1 : boolean;
  signal type_cast_2225_inst_ack_1 : boolean;
  signal phi_stmt_2222_req_0 : boolean;
  signal type_cast_2229_inst_req_0 : boolean;
  signal type_cast_2229_inst_ack_0 : boolean;
  signal type_cast_2229_inst_req_1 : boolean;
  signal type_cast_2229_inst_ack_1 : boolean;
  signal phi_stmt_2226_req_0 : boolean;
  signal phi_stmt_2218_ack_0 : boolean;
  signal phi_stmt_2222_ack_0 : boolean;
  signal phi_stmt_2226_ack_0 : boolean;
  signal type_cast_2337_inst_req_0 : boolean;
  signal type_cast_2337_inst_ack_0 : boolean;
  signal type_cast_2337_inst_req_1 : boolean;
  signal type_cast_2337_inst_ack_1 : boolean;
  signal phi_stmt_2331_req_1 : boolean;
  signal type_cast_2343_inst_req_0 : boolean;
  signal type_cast_2343_inst_ack_0 : boolean;
  signal type_cast_2343_inst_req_1 : boolean;
  signal type_cast_2343_inst_ack_1 : boolean;
  signal phi_stmt_2338_req_1 : boolean;
  signal type_cast_2349_inst_req_0 : boolean;
  signal type_cast_2349_inst_ack_0 : boolean;
  signal type_cast_2349_inst_req_1 : boolean;
  signal type_cast_2349_inst_ack_1 : boolean;
  signal phi_stmt_2344_req_1 : boolean;
  signal phi_stmt_2331_req_0 : boolean;
  signal type_cast_2341_inst_req_0 : boolean;
  signal type_cast_2341_inst_ack_0 : boolean;
  signal type_cast_2341_inst_req_1 : boolean;
  signal type_cast_2341_inst_ack_1 : boolean;
  signal phi_stmt_2338_req_0 : boolean;
  signal type_cast_2347_inst_req_0 : boolean;
  signal type_cast_2347_inst_ack_0 : boolean;
  signal type_cast_2347_inst_req_1 : boolean;
  signal type_cast_2347_inst_ack_1 : boolean;
  signal phi_stmt_2344_req_0 : boolean;
  signal phi_stmt_2331_ack_0 : boolean;
  signal phi_stmt_2338_ack_0 : boolean;
  signal phi_stmt_2344_ack_0 : boolean;
  signal phi_stmt_3397_req_0 : boolean;
  signal type_cast_3409_inst_req_0 : boolean;
  signal type_cast_3413_inst_ack_0 : boolean;
  signal phi_stmt_3410_req_1 : boolean;
  signal type_cast_3415_inst_ack_1 : boolean;
  signal type_cast_3415_inst_req_1 : boolean;
  signal type_cast_3415_inst_ack_0 : boolean;
  signal type_cast_3415_inst_req_0 : boolean;
  signal phi_stmt_2723_req_1 : boolean;
  signal type_cast_3413_inst_req_0 : boolean;
  signal type_cast_2735_inst_req_0 : boolean;
  signal type_cast_2735_inst_ack_0 : boolean;
  signal type_cast_2735_inst_req_1 : boolean;
  signal type_cast_2735_inst_ack_1 : boolean;
  signal phi_stmt_2730_req_1 : boolean;
  signal type_cast_2741_inst_req_0 : boolean;
  signal type_cast_2741_inst_ack_0 : boolean;
  signal type_cast_2741_inst_req_1 : boolean;
  signal type_cast_2741_inst_ack_1 : boolean;
  signal phi_stmt_2736_req_1 : boolean;
  signal type_cast_2726_inst_req_0 : boolean;
  signal type_cast_2726_inst_ack_0 : boolean;
  signal type_cast_2726_inst_req_1 : boolean;
  signal type_cast_2726_inst_ack_1 : boolean;
  signal phi_stmt_2723_req_0 : boolean;
  signal type_cast_2733_inst_req_0 : boolean;
  signal type_cast_2733_inst_ack_0 : boolean;
  signal type_cast_2733_inst_req_1 : boolean;
  signal type_cast_2733_inst_ack_1 : boolean;
  signal phi_stmt_2730_req_0 : boolean;
  signal phi_stmt_3814_req_1 : boolean;
  signal type_cast_2739_inst_req_0 : boolean;
  signal type_cast_2739_inst_ack_0 : boolean;
  signal type_cast_2739_inst_req_1 : boolean;
  signal type_cast_2739_inst_ack_1 : boolean;
  signal phi_stmt_2736_req_0 : boolean;
  signal type_cast_3819_inst_ack_1 : boolean;
  signal phi_stmt_2723_ack_0 : boolean;
  signal phi_stmt_2730_ack_0 : boolean;
  signal phi_stmt_2736_ack_0 : boolean;
  signal type_cast_3819_inst_req_1 : boolean;
  signal type_cast_2748_inst_req_0 : boolean;
  signal type_cast_2748_inst_ack_0 : boolean;
  signal type_cast_2748_inst_req_1 : boolean;
  signal type_cast_2748_inst_ack_1 : boolean;
  signal phi_stmt_3801_req_0 : boolean;
  signal phi_stmt_2745_req_0 : boolean;
  signal type_cast_3819_inst_ack_0 : boolean;
  signal type_cast_3819_inst_req_0 : boolean;
  signal type_cast_2752_inst_req_0 : boolean;
  signal type_cast_2752_inst_ack_0 : boolean;
  signal type_cast_2752_inst_req_1 : boolean;
  signal type_cast_2752_inst_ack_1 : boolean;
  signal phi_stmt_2749_req_0 : boolean;
  signal type_cast_3804_inst_ack_1 : boolean;
  signal phi_stmt_2745_ack_0 : boolean;
  signal phi_stmt_2749_ack_0 : boolean;
  signal type_cast_2850_inst_req_0 : boolean;
  signal type_cast_2850_inst_ack_0 : boolean;
  signal type_cast_2850_inst_req_1 : boolean;
  signal phi_stmt_3410_ack_0 : boolean;
  signal type_cast_2850_inst_ack_1 : boolean;
  signal type_cast_3804_inst_req_1 : boolean;
  signal phi_stmt_2844_req_1 : boolean;
  signal type_cast_2856_inst_req_0 : boolean;
  signal type_cast_2856_inst_ack_0 : boolean;
  signal phi_stmt_3404_ack_0 : boolean;
  signal type_cast_2856_inst_req_1 : boolean;
  signal phi_stmt_3397_ack_0 : boolean;
  signal type_cast_2856_inst_ack_1 : boolean;
  signal phi_stmt_2851_req_1 : boolean;
  signal phi_stmt_3404_req_0 : boolean;
  signal type_cast_2863_inst_req_0 : boolean;
  signal type_cast_2863_inst_ack_0 : boolean;
  signal type_cast_2863_inst_req_1 : boolean;
  signal type_cast_2863_inst_ack_1 : boolean;
  signal phi_stmt_2857_req_1 : boolean;
  signal phi_stmt_3410_req_0 : boolean;
  signal phi_stmt_2844_req_0 : boolean;
  signal phi_stmt_3404_req_1 : boolean;
  signal type_cast_2854_inst_req_0 : boolean;
  signal type_cast_2854_inst_ack_0 : boolean;
  signal type_cast_3413_inst_ack_1 : boolean;
  signal type_cast_2854_inst_req_1 : boolean;
  signal type_cast_2854_inst_ack_1 : boolean;
  signal phi_stmt_2851_req_0 : boolean;
  signal phi_stmt_2857_req_0 : boolean;
  signal type_cast_3413_inst_req_1 : boolean;
  signal type_cast_3407_inst_ack_1 : boolean;
  signal phi_stmt_2844_ack_0 : boolean;
  signal phi_stmt_2851_ack_0 : boolean;
  signal phi_stmt_2857_ack_0 : boolean;
  signal type_cast_3278_inst_req_0 : boolean;
  signal type_cast_3278_inst_ack_0 : boolean;
  signal type_cast_3278_inst_req_1 : boolean;
  signal type_cast_3278_inst_ack_1 : boolean;
  signal phi_stmt_3275_req_0 : boolean;
  signal type_cast_3274_inst_req_0 : boolean;
  signal type_cast_3274_inst_ack_0 : boolean;
  signal type_cast_3274_inst_req_1 : boolean;
  signal type_cast_3274_inst_ack_1 : boolean;
  signal phi_stmt_3269_req_1 : boolean;
  signal phi_stmt_3262_req_0 : boolean;
  signal type_cast_3280_inst_req_0 : boolean;
  signal type_cast_3280_inst_ack_0 : boolean;
  signal type_cast_3280_inst_req_1 : boolean;
  signal type_cast_3280_inst_ack_1 : boolean;
  signal phi_stmt_3275_req_1 : boolean;
  signal type_cast_3272_inst_req_0 : boolean;
  signal type_cast_3272_inst_ack_0 : boolean;
  signal type_cast_3272_inst_req_1 : boolean;
  signal type_cast_3272_inst_ack_1 : boolean;
  signal phi_stmt_3269_req_0 : boolean;
  signal type_cast_3268_inst_req_0 : boolean;
  signal type_cast_3268_inst_ack_0 : boolean;
  signal type_cast_3268_inst_req_1 : boolean;
  signal type_cast_3268_inst_ack_1 : boolean;
  signal phi_stmt_3262_req_1 : boolean;
  signal phi_stmt_3262_ack_0 : boolean;
  signal phi_stmt_3269_ack_0 : boolean;
  signal phi_stmt_3275_ack_0 : boolean;
  signal type_cast_3295_inst_req_0 : boolean;
  signal type_cast_3295_inst_ack_0 : boolean;
  signal type_cast_3295_inst_req_1 : boolean;
  signal type_cast_3295_inst_ack_1 : boolean;
  signal phi_stmt_3292_req_0 : boolean;
  signal type_cast_3291_inst_req_0 : boolean;
  signal type_cast_3291_inst_ack_0 : boolean;
  signal type_cast_3291_inst_req_1 : boolean;
  signal type_cast_3291_inst_ack_1 : boolean;
  signal phi_stmt_3288_req_0 : boolean;
  signal type_cast_3287_inst_req_0 : boolean;
  signal type_cast_3287_inst_ack_0 : boolean;
  signal type_cast_3287_inst_req_1 : boolean;
  signal type_cast_3287_inst_ack_1 : boolean;
  signal phi_stmt_3284_req_0 : boolean;
  signal phi_stmt_3284_ack_0 : boolean;
  signal phi_stmt_3288_ack_0 : boolean;
  signal phi_stmt_3292_ack_0 : boolean;
  signal type_cast_3403_inst_req_0 : boolean;
  signal type_cast_3403_inst_ack_0 : boolean;
  signal type_cast_3403_inst_req_1 : boolean;
  signal type_cast_3403_inst_ack_1 : boolean;
  signal phi_stmt_3397_req_1 : boolean;
  signal type_cast_3407_inst_req_0 : boolean;
  signal type_cast_3407_inst_ack_0 : boolean;
  signal type_cast_3407_inst_req_1 : boolean;
  signal type_cast_3811_inst_req_0 : boolean;
  signal type_cast_3811_inst_ack_0 : boolean;
  signal type_cast_3811_inst_req_1 : boolean;
  signal type_cast_3811_inst_ack_1 : boolean;
  signal phi_stmt_3808_req_0 : boolean;
  signal type_cast_3817_inst_req_0 : boolean;
  signal type_cast_3817_inst_ack_0 : boolean;
  signal type_cast_3817_inst_req_1 : boolean;
  signal type_cast_3817_inst_ack_1 : boolean;
  signal phi_stmt_3814_req_0 : boolean;
  signal phi_stmt_3801_ack_0 : boolean;
  signal phi_stmt_3808_ack_0 : boolean;
  signal phi_stmt_3814_ack_0 : boolean;
  signal type_cast_3826_inst_req_0 : boolean;
  signal type_cast_3826_inst_ack_0 : boolean;
  signal type_cast_3826_inst_req_1 : boolean;
  signal type_cast_3826_inst_ack_1 : boolean;
  signal phi_stmt_3823_req_0 : boolean;
  signal type_cast_3830_inst_req_0 : boolean;
  signal type_cast_3830_inst_ack_0 : boolean;
  signal type_cast_3830_inst_req_1 : boolean;
  signal type_cast_3830_inst_ack_1 : boolean;
  signal phi_stmt_3827_req_0 : boolean;
  signal phi_stmt_3823_ack_0 : boolean;
  signal phi_stmt_3827_ack_0 : boolean;
  signal type_cast_3934_inst_req_0 : boolean;
  signal type_cast_3934_inst_ack_0 : boolean;
  signal type_cast_3934_inst_req_1 : boolean;
  signal type_cast_3934_inst_ack_1 : boolean;
  signal phi_stmt_3928_req_1 : boolean;
  signal type_cast_3938_inst_req_0 : boolean;
  signal type_cast_3938_inst_ack_0 : boolean;
  signal type_cast_3938_inst_req_1 : boolean;
  signal type_cast_3938_inst_ack_1 : boolean;
  signal phi_stmt_3935_req_0 : boolean;
  signal type_cast_3947_inst_req_0 : boolean;
  signal type_cast_3947_inst_ack_0 : boolean;
  signal type_cast_3947_inst_req_1 : boolean;
  signal type_cast_3947_inst_ack_1 : boolean;
  signal phi_stmt_3941_req_1 : boolean;
  signal phi_stmt_3928_req_0 : boolean;
  signal type_cast_3940_inst_req_0 : boolean;
  signal type_cast_3940_inst_ack_0 : boolean;
  signal type_cast_3940_inst_req_1 : boolean;
  signal type_cast_3940_inst_ack_1 : boolean;
  signal phi_stmt_3935_req_1 : boolean;
  signal phi_stmt_3941_req_0 : boolean;
  signal phi_stmt_3928_ack_0 : boolean;
  signal phi_stmt_3935_ack_0 : boolean;
  signal phi_stmt_3941_ack_0 : boolean;
  signal phi_stmt_4322_req_1 : boolean;
  signal type_cast_4334_inst_req_0 : boolean;
  signal type_cast_4334_inst_ack_0 : boolean;
  signal type_cast_4334_inst_req_1 : boolean;
  signal type_cast_4334_inst_ack_1 : boolean;
  signal phi_stmt_4329_req_1 : boolean;
  signal type_cast_4340_inst_req_0 : boolean;
  signal type_cast_4340_inst_ack_0 : boolean;
  signal type_cast_4340_inst_req_1 : boolean;
  signal type_cast_4340_inst_ack_1 : boolean;
  signal phi_stmt_4335_req_1 : boolean;
  signal type_cast_4325_inst_req_0 : boolean;
  signal type_cast_4325_inst_ack_0 : boolean;
  signal type_cast_4325_inst_req_1 : boolean;
  signal type_cast_4325_inst_ack_1 : boolean;
  signal phi_stmt_4322_req_0 : boolean;
  signal type_cast_4332_inst_req_0 : boolean;
  signal type_cast_4332_inst_ack_0 : boolean;
  signal type_cast_4332_inst_req_1 : boolean;
  signal type_cast_4332_inst_ack_1 : boolean;
  signal phi_stmt_4329_req_0 : boolean;
  signal type_cast_4338_inst_req_0 : boolean;
  signal type_cast_4338_inst_ack_0 : boolean;
  signal type_cast_4338_inst_req_1 : boolean;
  signal type_cast_4338_inst_ack_1 : boolean;
  signal phi_stmt_4335_req_0 : boolean;
  signal phi_stmt_4322_ack_0 : boolean;
  signal phi_stmt_4329_ack_0 : boolean;
  signal phi_stmt_4335_ack_0 : boolean;
  signal type_cast_4347_inst_req_0 : boolean;
  signal type_cast_4347_inst_ack_0 : boolean;
  signal type_cast_4347_inst_req_1 : boolean;
  signal type_cast_4347_inst_ack_1 : boolean;
  signal phi_stmt_4344_req_0 : boolean;
  signal type_cast_4351_inst_req_0 : boolean;
  signal type_cast_4351_inst_ack_0 : boolean;
  signal type_cast_4351_inst_req_1 : boolean;
  signal type_cast_4351_inst_ack_1 : boolean;
  signal phi_stmt_4348_req_0 : boolean;
  signal type_cast_4355_inst_req_0 : boolean;
  signal type_cast_4355_inst_ack_0 : boolean;
  signal type_cast_4355_inst_req_1 : boolean;
  signal type_cast_4355_inst_ack_1 : boolean;
  signal phi_stmt_4352_req_0 : boolean;
  signal phi_stmt_4344_ack_0 : boolean;
  signal phi_stmt_4348_ack_0 : boolean;
  signal phi_stmt_4352_ack_0 : boolean;
  signal type_cast_4469_inst_req_0 : boolean;
  signal type_cast_4469_inst_ack_0 : boolean;
  signal type_cast_4469_inst_req_1 : boolean;
  signal type_cast_4469_inst_ack_1 : boolean;
  signal phi_stmt_4463_req_1 : boolean;
  signal type_cast_4475_inst_req_0 : boolean;
  signal type_cast_4475_inst_ack_0 : boolean;
  signal type_cast_4475_inst_req_1 : boolean;
  signal type_cast_4475_inst_ack_1 : boolean;
  signal phi_stmt_4470_req_1 : boolean;
  signal type_cast_4481_inst_req_0 : boolean;
  signal type_cast_4481_inst_ack_0 : boolean;
  signal type_cast_4481_inst_req_1 : boolean;
  signal type_cast_4481_inst_ack_1 : boolean;
  signal phi_stmt_4476_req_1 : boolean;
  signal phi_stmt_4463_req_0 : boolean;
  signal type_cast_4473_inst_req_0 : boolean;
  signal type_cast_4473_inst_ack_0 : boolean;
  signal type_cast_4473_inst_req_1 : boolean;
  signal type_cast_4473_inst_ack_1 : boolean;
  signal phi_stmt_4470_req_0 : boolean;
  signal type_cast_4479_inst_req_0 : boolean;
  signal type_cast_4479_inst_ack_0 : boolean;
  signal type_cast_4479_inst_req_1 : boolean;
  signal type_cast_4479_inst_ack_1 : boolean;
  signal phi_stmt_4476_req_0 : boolean;
  signal phi_stmt_4463_ack_0 : boolean;
  signal phi_stmt_4470_ack_0 : boolean;
  signal phi_stmt_4476_ack_0 : boolean;
  signal type_cast_4861_inst_req_0 : boolean;
  signal type_cast_4861_inst_ack_0 : boolean;
  signal type_cast_4861_inst_req_1 : boolean;
  signal type_cast_4861_inst_ack_1 : boolean;
  signal phi_stmt_4856_req_1 : boolean;
  signal phi_stmt_4843_req_0 : boolean;
  signal type_cast_4855_inst_req_0 : boolean;
  signal type_cast_4855_inst_ack_0 : boolean;
  signal type_cast_4855_inst_req_1 : boolean;
  signal type_cast_4855_inst_ack_1 : boolean;
  signal phi_stmt_4850_req_1 : boolean;
  signal type_cast_4859_inst_req_0 : boolean;
  signal type_cast_4859_inst_ack_0 : boolean;
  signal type_cast_4859_inst_req_1 : boolean;
  signal type_cast_4859_inst_ack_1 : boolean;
  signal phi_stmt_4856_req_0 : boolean;
  signal type_cast_4849_inst_req_0 : boolean;
  signal type_cast_4849_inst_ack_0 : boolean;
  signal type_cast_4849_inst_req_1 : boolean;
  signal type_cast_4849_inst_ack_1 : boolean;
  signal phi_stmt_4843_req_1 : boolean;
  signal type_cast_4853_inst_req_0 : boolean;
  signal type_cast_4853_inst_ack_0 : boolean;
  signal type_cast_4853_inst_req_1 : boolean;
  signal type_cast_4853_inst_ack_1 : boolean;
  signal phi_stmt_4850_req_0 : boolean;
  signal phi_stmt_4843_ack_0 : boolean;
  signal phi_stmt_4850_ack_0 : boolean;
  signal phi_stmt_4856_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_2067_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2067_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_2067_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2067_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_2067: Block -- control-path 
    signal zeropad3D_CP_2067_elements: BooleanArray(1250 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_2067_elements(0) <= zeropad3D_CP_2067_start;
    zeropad3D_CP_2067_symbol <= zeropad3D_CP_2067_elements(796);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_update_start_
      -- CP-element group 0: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_655/call_stmt_657/$entry
      -- CP-element group 0: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_Update/ccr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_655/$entry
      -- CP-element group 0: 	 branch_block_stmt_655/branch_block_stmt_655__entry__
      -- CP-element group 0: 	 branch_block_stmt_655/call_stmt_657__entry__
      -- 
    crr_2523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(0), ack => call_stmt_657_call_req_0); -- 
    ccr_2528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(0), ack => call_stmt_657_call_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	840 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	801 
    -- CP-element group 1: 	802 
    -- CP-element group 1: 	804 
    -- CP-element group 1: 	805 
    -- CP-element group 1: 	807 
    -- CP-element group 1: 	808 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_655/merge_stmt_1154__exit__
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/Update/cr
      -- 
    rr_10699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1), ack => type_cast_753_inst_req_0); -- 
    cr_10704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1), ack => type_cast_753_inst_req_1); -- 
    rr_10722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1), ack => type_cast_760_inst_req_0); -- 
    cr_10727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1), ack => type_cast_760_inst_req_1); -- 
    rr_10745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1), ack => type_cast_767_inst_req_0); -- 
    cr_10750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1), ack => type_cast_767_inst_req_1); -- 
    zeropad3D_CP_2067_elements(1) <= zeropad3D_CP_2067_elements(840);
    -- CP-element group 2:  merge  fork  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	896 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	851 
    -- CP-element group 2: 	852 
    -- CP-element group 2: 	854 
    -- CP-element group 2: 	855 
    -- CP-element group 2: 	857 
    -- CP-element group 2: 	858 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_655/merge_stmt_1668__exit__
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Update/cr
      -- 
    rr_11069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(2), ack => type_cast_1281_inst_req_0); -- 
    cr_11074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(2), ack => type_cast_1281_inst_req_1); -- 
    rr_11092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(2), ack => type_cast_1288_inst_req_0); -- 
    cr_11097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(2), ack => type_cast_1288_inst_req_1); -- 
    rr_11115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(2), ack => type_cast_1295_inst_req_0); -- 
    cr_11120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(2), ack => type_cast_1295_inst_req_1); -- 
    zeropad3D_CP_2067_elements(2) <= zeropad3D_CP_2067_elements(896);
    -- CP-element group 3:  merge  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	952 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	907 
    -- CP-element group 3: 	908 
    -- CP-element group 3: 	910 
    -- CP-element group 3: 	911 
    -- CP-element group 3: 	913 
    -- CP-element group 3: 	914 
    -- CP-element group 3:  members (27) 
      -- CP-element group 3: 	 branch_block_stmt_655/merge_stmt_2195__exit__
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/$entry
      -- CP-element group 3: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Sample/$entry
      -- 
    rr_11481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(3), ack => type_cast_1809_inst_req_0); -- 
    cr_11532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(3), ack => type_cast_1793_inst_req_1); -- 
    rr_11527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(3), ack => type_cast_1793_inst_req_0); -- 
    cr_11486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(3), ack => type_cast_1809_inst_req_1); -- 
    cr_11509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(3), ack => type_cast_1802_inst_req_1); -- 
    rr_11504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(3), ack => type_cast_1802_inst_req_0); -- 
    zeropad3D_CP_2067_elements(3) <= zeropad3D_CP_2067_elements(952);
    -- CP-element group 4:  merge  fork  transition  place  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1014 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	967 
    -- CP-element group 4: 	968 
    -- CP-element group 4: 	970 
    -- CP-element group 4: 	971 
    -- CP-element group 4: 	973 
    -- CP-element group 4: 	974 
    -- CP-element group 4:  members (27) 
      -- CP-element group 4: 	 branch_block_stmt_655/merge_stmt_2722__exit__
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/Update/cr
      -- 
    rr_11917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(4), ack => type_cast_2337_inst_req_0); -- 
    cr_11922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(4), ack => type_cast_2337_inst_req_1); -- 
    rr_11940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(4), ack => type_cast_2343_inst_req_0); -- 
    cr_11945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(4), ack => type_cast_2343_inst_req_1); -- 
    rr_11963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(4), ack => type_cast_2349_inst_req_0); -- 
    cr_11968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(4), ack => type_cast_2349_inst_req_1); -- 
    zeropad3D_CP_2067_elements(4) <= zeropad3D_CP_2067_elements(1014);
    -- CP-element group 5:  merge  fork  transition  place  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1070 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	1025 
    -- CP-element group 5: 	1026 
    -- CP-element group 5: 	1028 
    -- CP-element group 5: 	1029 
    -- CP-element group 5: 	1031 
    -- CP-element group 5: 	1032 
    -- CP-element group 5:  members (27) 
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888
      -- CP-element group 5: 	 branch_block_stmt_655/merge_stmt_3261__exit__
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/Update/cr
      -- 
    rr_12344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(5), ack => type_cast_2850_inst_req_0); -- 
    cr_12349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(5), ack => type_cast_2850_inst_req_1); -- 
    rr_12367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(5), ack => type_cast_2856_inst_req_0); -- 
    cr_12372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(5), ack => type_cast_2856_inst_req_1); -- 
    rr_12390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(5), ack => type_cast_2863_inst_req_0); -- 
    cr_12395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(5), ack => type_cast_2863_inst_req_1); -- 
    zeropad3D_CP_2067_elements(5) <= zeropad3D_CP_2067_elements(1070);
    -- CP-element group 6:  merge  fork  transition  place  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1132 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	1085 
    -- CP-element group 6: 	1086 
    -- CP-element group 6: 	1088 
    -- CP-element group 6: 	1089 
    -- CP-element group 6: 	1091 
    -- CP-element group 6: 	1092 
    -- CP-element group 6:  members (27) 
      -- CP-element group 6: 	 branch_block_stmt_655/merge_stmt_3800__exit__
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/Update/cr
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/Update/cr
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/Update/cr
      -- 
    cr_12831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(6), ack => type_cast_3415_inst_req_1); -- 
    rr_12826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(6), ack => type_cast_3415_inst_req_0); -- 
    rr_12780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(6), ack => type_cast_3403_inst_req_0); -- 
    cr_12785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(6), ack => type_cast_3403_inst_req_1); -- 
    rr_12803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(6), ack => type_cast_3407_inst_req_0); -- 
    cr_12808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(6), ack => type_cast_3407_inst_req_1); -- 
    zeropad3D_CP_2067_elements(6) <= zeropad3D_CP_2067_elements(1132);
    -- CP-element group 7:  merge  fork  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1188 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	1143 
    -- CP-element group 7: 	1144 
    -- CP-element group 7: 	1146 
    -- CP-element group 7: 	1147 
    -- CP-element group 7: 	1149 
    -- CP-element group 7: 	1150 
    -- CP-element group 7:  members (27) 
      -- CP-element group 7: 	 branch_block_stmt_655/merge_stmt_4321__exit__
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/Update/cr
      -- 
    rr_13207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(7), ack => type_cast_3934_inst_req_0); -- 
    cr_13212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(7), ack => type_cast_3934_inst_req_1); -- 
    rr_13230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(7), ack => type_cast_3938_inst_req_0); -- 
    cr_13235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(7), ack => type_cast_3938_inst_req_1); -- 
    rr_13253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(7), ack => type_cast_3947_inst_req_0); -- 
    cr_13258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(7), ack => type_cast_3947_inst_req_1); -- 
    zeropad3D_CP_2067_elements(7) <= zeropad3D_CP_2067_elements(1188);
    -- CP-element group 8:  merge  fork  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1250 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	1203 
    -- CP-element group 8: 	1204 
    -- CP-element group 8: 	1206 
    -- CP-element group 8: 	1207 
    -- CP-element group 8: 	1209 
    -- CP-element group 8: 	1210 
    -- CP-element group 8:  members (27) 
      -- CP-element group 8: 	 branch_block_stmt_655/merge_stmt_4842__exit__
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/Update/cr
      -- 
    rr_13643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(8), ack => type_cast_4469_inst_req_0); -- 
    cr_13648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(8), ack => type_cast_4469_inst_req_1); -- 
    rr_13666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(8), ack => type_cast_4475_inst_req_0); -- 
    cr_13671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(8), ack => type_cast_4475_inst_req_1); -- 
    rr_13689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(8), ack => type_cast_4481_inst_req_0); -- 
    cr_13694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(8), ack => type_cast_4481_inst_req_1); -- 
    zeropad3D_CP_2067_elements(8) <= zeropad3D_CP_2067_elements(1250);
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_Sample/cra
      -- 
    cra_2524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_657_call_ack_0, ack => zeropad3D_CP_2067_elements(9)); -- 
    -- CP-element group 10:  fork  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	18 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	20 
    -- CP-element group 10: 	22 
    -- CP-element group 10: 	24 
    -- CP-element group 10: 	26 
    -- CP-element group 10: 	28 
    -- CP-element group 10: 	30 
    -- CP-element group 10: 	32 
    -- CP-element group 10:  members (85) 
      -- CP-element group 10: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_Update/cca
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/word_access_complete/word_0/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Sample/word_access_start/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/word_access_complete/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/word_access_complete/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Sample/word_access_start/word_0/rr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Sample/word_access_start/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Sample/word_access_start/word_0/rr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Sample/word_access_start/word_0/rr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/word_access_complete/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Sample/word_access_start/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/word_access_complete/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/word_access_complete/word_0/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_word_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_root_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Sample/word_access_start/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_word_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/word_access_complete/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/word_access_complete/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_root_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Sample/word_access_start/word_0/rr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Sample/word_access_start/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Sample/word_access_start/word_0/rr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_word_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/call_stmt_657/call_stmt_657_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_root_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/word_access_complete/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_word_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/word_access_complete/word_0/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_root_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/call_stmt_657/$exit
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/word_access_complete/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/word_access_complete/word_0/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_root_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_word_address_calculated
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/word_access_complete/word_0/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/word_access_complete/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/word_access_complete/word_0/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/call_stmt_657__exit__
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744__entry__
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_update_start_
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_Update/cr
      -- 
    cca_2529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_657_call_ack_1, ack => zeropad3D_CP_2067_elements(10)); -- 
    cr_2559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_pad_660_load_0_req_1); -- 
    rr_2548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_pad_660_load_0_req_0); -- 
    rr_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_out_depth_high_669_load_0_req_0); -- 
    rr_2581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_depth_high_663_load_0_req_0); -- 
    cr_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_depth_high_663_load_0_req_1); -- 
    rr_2614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_col_high_666_load_0_req_0); -- 
    rr_2680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_out_col_high_672_load_0_req_0); -- 
    cr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_out_depth_high_669_load_0_req_1); -- 
    cr_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_col_high_666_load_0_req_1); -- 
    cr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => LOAD_out_col_high_672_load_0_req_1); -- 
    cr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => type_cast_676_inst_req_1); -- 
    cr_2724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => type_cast_680_inst_req_1); -- 
    cr_2738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => type_cast_684_inst_req_1); -- 
    cr_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => type_cast_688_inst_req_1); -- 
    cr_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => type_cast_697_inst_req_1); -- 
    cr_2780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(10), ack => type_cast_701_inst_req_1); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Sample/word_access_start/word_0/ra
      -- 
    ra_2549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_660_load_0_ack_0, ack => zeropad3D_CP_2067_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (12) 
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/LOAD_pad_660_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/LOAD_pad_660_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/LOAD_pad_660_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_pad_660_Update/LOAD_pad_660_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_Sample/rr
      -- 
    ca_2560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_660_load_0_ack_1, ack => zeropad3D_CP_2067_elements(12)); -- 
    rr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(12), ack => type_cast_697_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Sample/$exit
      -- 
    ra_2582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_663_load_0_ack_0, ack => zeropad3D_CP_2067_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	21 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/LOAD_depth_high_663_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/LOAD_depth_high_663_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/LOAD_depth_high_663_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_Update/LOAD_depth_high_663_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_depth_high_663_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_Sample/rr
      -- 
    ca_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_663_load_0_ack_1, ack => zeropad3D_CP_2067_elements(14)); -- 
    rr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(14), ack => type_cast_676_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Sample/word_access_start/word_0/$exit
      -- 
    ra_2615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_666_load_0_ack_0, ack => zeropad3D_CP_2067_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	23 
    -- CP-element group 16:  members (12) 
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/LOAD_col_high_666_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/LOAD_col_high_666_Merge/merge_ack
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/LOAD_col_high_666_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/LOAD_col_high_666_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_col_high_666_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_Sample/rr
      -- 
    ca_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_666_load_0_ack_1, ack => zeropad3D_CP_2067_elements(16)); -- 
    rr_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(16), ack => type_cast_680_inst_req_0); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Sample/word_access_start/word_0/ra
      -- CP-element group 17: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Sample/word_access_start/$exit
      -- 
    ra_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_669_load_0_ack_0, ack => zeropad3D_CP_2067_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	10 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	31 
    -- CP-element group 18:  members (15) 
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/LOAD_out_depth_high_669_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/LOAD_out_depth_high_669_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/LOAD_out_depth_high_669_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_depth_high_669_Update/LOAD_out_depth_high_669_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_Sample/rr
      -- 
    ca_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_669_load_0_ack_1, ack => zeropad3D_CP_2067_elements(18)); -- 
    rr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(18), ack => type_cast_684_inst_req_0); -- 
    rr_2775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(18), ack => type_cast_701_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Sample/$exit
      -- 
    ra_2681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_672_load_0_ack_0, ack => zeropad3D_CP_2067_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	27 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/LOAD_out_col_high_672_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/LOAD_out_col_high_672_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/LOAD_out_col_high_672_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/LOAD_out_col_high_672_Update/LOAD_out_col_high_672_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_Sample/rr
      -- 
    ca_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_672_load_0_ack_1, ack => zeropad3D_CP_2067_elements(20)); -- 
    rr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(20), ack => type_cast_688_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_Sample/ra
      -- 
    ra_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_676_inst_ack_0, ack => zeropad3D_CP_2067_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	10 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	33 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_676_Update/ca
      -- 
    ca_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_676_inst_ack_1, ack => zeropad3D_CP_2067_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_Sample/ra
      -- 
    ra_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_680_inst_ack_0, ack => zeropad3D_CP_2067_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	10 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	33 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_680_Update/ca
      -- 
    ca_2725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_680_inst_ack_1, ack => zeropad3D_CP_2067_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_Sample/ra
      -- 
    ra_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_684_inst_ack_0, ack => zeropad3D_CP_2067_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	10 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	33 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_684_Update/ca
      -- 
    ca_2739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_684_inst_ack_1, ack => zeropad3D_CP_2067_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	20 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_Sample/ra
      -- 
    ra_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_0, ack => zeropad3D_CP_2067_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	10 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	33 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_688_Update/ca
      -- 
    ca_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_1, ack => zeropad3D_CP_2067_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	12 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_Sample/ra
      -- 
    ra_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_697_inst_ack_0, ack => zeropad3D_CP_2067_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	10 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_697_Update/ca
      -- 
    ca_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_697_inst_ack_1, ack => zeropad3D_CP_2067_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	18 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_Sample/ra
      -- 
    ra_2776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_0, ack => zeropad3D_CP_2067_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	10 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/type_cast_701_Update/ca
      -- 
    ca_2781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_1, ack => zeropad3D_CP_2067_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  place  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	24 
    -- CP-element group 33: 	26 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	30 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	797 
    -- CP-element group 33: 	798 
    -- CP-element group 33: 	799 
    -- CP-element group 33:  members (10) 
      -- CP-element group 33: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744/$exit
      -- CP-element group 33: 	 branch_block_stmt_655/assign_stmt_661_to_assign_stmt_744__exit__
      -- CP-element group 33: 	 branch_block_stmt_655/entry_whilex_xbody
      -- CP-element group 33: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_747/$entry
      -- CP-element group 33: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_754/$entry
      -- CP-element group 33: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_761/$entry
      -- CP-element group 33: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/$entry
      -- 
    zeropad3D_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(22) & zeropad3D_CP_2067_elements(24) & zeropad3D_CP_2067_elements(26) & zeropad3D_CP_2067_elements(28) & zeropad3D_CP_2067_elements(30) & zeropad3D_CP_2067_elements(32);
      gj_zeropad3D_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	815 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_Sample/ra
      -- 
    ra_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_772_inst_ack_0, ack => zeropad3D_CP_2067_elements(34)); -- 
    -- CP-element group 35:  branch  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	815 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (13) 
      -- CP-element group 35: 	 branch_block_stmt_655/R_cmp_782_place
      -- CP-element group 35: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780__exit__
      -- CP-element group 35: 	 branch_block_stmt_655/if_stmt_781__entry__
      -- CP-element group 35: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/$exit
      -- CP-element group 35: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_655/if_stmt_781_dead_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_655/if_stmt_781_eval_test/$entry
      -- CP-element group 35: 	 branch_block_stmt_655/if_stmt_781_eval_test/$exit
      -- CP-element group 35: 	 branch_block_stmt_655/if_stmt_781_eval_test/branch_req
      -- CP-element group 35: 	 branch_block_stmt_655/if_stmt_781_if_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_655/if_stmt_781_else_link/$entry
      -- 
    ca_2798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_772_inst_ack_1, ack => zeropad3D_CP_2067_elements(35)); -- 
    branch_req_2806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(35), ack => if_stmt_781_branch_req_0); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	816 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_655/whilex_xbody_ifx_xthen
      -- CP-element group 36: 	 branch_block_stmt_655/if_stmt_781_if_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_655/if_stmt_781_if_link/if_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_655/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_655/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    if_choice_transition_2811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_781_branch_ack_1, ack => zeropad3D_CP_2067_elements(36)); -- 
    -- CP-element group 37:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	41 
    -- CP-element group 37:  members (27) 
      -- CP-element group 37: 	 branch_block_stmt_655/merge_stmt_787__exit__
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812__entry__
      -- CP-element group 37: 	 branch_block_stmt_655/if_stmt_781_else_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_655/if_stmt_781_else_link/else_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_655/whilex_xbody_lorx_xlhsx_xfalse
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_update_start_
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_word_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Sample/word_access_start/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Sample/word_access_start/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Sample/word_access_start/word_0/rr
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/word_access_complete/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/word_access_complete/word_0/cr
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_update_start_
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_655/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_655/merge_stmt_787_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_655/merge_stmt_787_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_655/merge_stmt_787_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_655/merge_stmt_787_PhiAck/dummy
      -- 
    else_choice_transition_2815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_781_branch_ack_0, ack => zeropad3D_CP_2067_elements(37)); -- 
    rr_2836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(37), ack => LOAD_row_high_789_load_0_req_0); -- 
    cr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(37), ack => LOAD_row_high_789_load_0_req_1); -- 
    cr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(37), ack => type_cast_793_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Sample/word_access_start/$exit
      -- CP-element group 38: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Sample/word_access_start/word_0/ra
      -- 
    ra_2837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_789_load_0_ack_0, ack => zeropad3D_CP_2067_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (12) 
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/word_access_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/LOAD_row_high_789_Merge/$entry
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/LOAD_row_high_789_Merge/$exit
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/LOAD_row_high_789_Merge/merge_req
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/LOAD_row_high_789_Update/LOAD_row_high_789_Merge/merge_ack
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_Sample/rr
      -- 
    ca_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_789_load_0_ack_1, ack => zeropad3D_CP_2067_elements(39)); -- 
    rr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(39), ack => type_cast_793_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_Sample/ra
      -- 
    ra_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_0, ack => zeropad3D_CP_2067_elements(40)); -- 
    -- CP-element group 41:  branch  transition  place  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	37 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (13) 
      -- CP-element group 41: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812__exit__
      -- CP-element group 41: 	 branch_block_stmt_655/if_stmt_813__entry__
      -- CP-element group 41: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/$exit
      -- CP-element group 41: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_655/assign_stmt_790_to_assign_stmt_812/type_cast_793_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_655/if_stmt_813_dead_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_655/if_stmt_813_eval_test/$entry
      -- CP-element group 41: 	 branch_block_stmt_655/if_stmt_813_eval_test/$exit
      -- CP-element group 41: 	 branch_block_stmt_655/if_stmt_813_eval_test/branch_req
      -- CP-element group 41: 	 branch_block_stmt_655/R_cmp46_814_place
      -- CP-element group 41: 	 branch_block_stmt_655/if_stmt_813_if_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_655/if_stmt_813_else_link/$entry
      -- 
    ca_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_1, ack => zeropad3D_CP_2067_elements(41)); -- 
    branch_req_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(41), ack => if_stmt_813_branch_req_0); -- 
    -- CP-element group 42:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (18) 
      -- CP-element group 42: 	 branch_block_stmt_655/merge_stmt_819__exit__
      -- CP-element group 42: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831__entry__
      -- CP-element group 42: 	 branch_block_stmt_655/if_stmt_813_if_link/$exit
      -- CP-element group 42: 	 branch_block_stmt_655/if_stmt_813_if_link/if_choice_transition
      -- CP-element group 42: 	 branch_block_stmt_655/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse48
      -- CP-element group 42: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/$entry
      -- CP-element group 42: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_update_start_
      -- CP-element group 42: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_Update/cr
      -- CP-element group 42: 	 branch_block_stmt_655/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse48_PhiReq/$entry
      -- CP-element group 42: 	 branch_block_stmt_655/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse48_PhiReq/$exit
      -- CP-element group 42: 	 branch_block_stmt_655/merge_stmt_819_PhiReqMerge
      -- CP-element group 42: 	 branch_block_stmt_655/merge_stmt_819_PhiAck/$entry
      -- CP-element group 42: 	 branch_block_stmt_655/merge_stmt_819_PhiAck/$exit
      -- CP-element group 42: 	 branch_block_stmt_655/merge_stmt_819_PhiAck/dummy
      -- 
    if_choice_transition_2880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_813_branch_ack_1, ack => zeropad3D_CP_2067_elements(42)); -- 
    rr_2897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(42), ack => type_cast_823_inst_req_0); -- 
    cr_2902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(42), ack => type_cast_823_inst_req_1); -- 
    -- CP-element group 43:  transition  place  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	816 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_655/if_stmt_813_else_link/$exit
      -- CP-element group 43: 	 branch_block_stmt_655/if_stmt_813_else_link/else_choice_transition
      -- CP-element group 43: 	 branch_block_stmt_655/lorx_xlhsx_xfalse_ifx_xthen
      -- CP-element group 43: 	 branch_block_stmt_655/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_655/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_2884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_813_branch_ack_0, ack => zeropad3D_CP_2067_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_Sample/ra
      -- 
    ra_2898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_0, ack => zeropad3D_CP_2067_elements(44)); -- 
    -- CP-element group 45:  branch  transition  place  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (13) 
      -- CP-element group 45: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831__exit__
      -- CP-element group 45: 	 branch_block_stmt_655/if_stmt_832__entry__
      -- CP-element group 45: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/$exit
      -- CP-element group 45: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_655/assign_stmt_824_to_assign_stmt_831/type_cast_823_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_655/if_stmt_832_dead_link/$entry
      -- CP-element group 45: 	 branch_block_stmt_655/if_stmt_832_eval_test/$entry
      -- CP-element group 45: 	 branch_block_stmt_655/if_stmt_832_eval_test/$exit
      -- CP-element group 45: 	 branch_block_stmt_655/if_stmt_832_eval_test/branch_req
      -- CP-element group 45: 	 branch_block_stmt_655/R_cmp53_833_place
      -- CP-element group 45: 	 branch_block_stmt_655/if_stmt_832_if_link/$entry
      -- CP-element group 45: 	 branch_block_stmt_655/if_stmt_832_else_link/$entry
      -- 
    ca_2903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_1, ack => zeropad3D_CP_2067_elements(45)); -- 
    branch_req_2911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(45), ack => if_stmt_832_branch_req_0); -- 
    -- CP-element group 46:  transition  place  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	816 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_655/if_stmt_832_if_link/$exit
      -- CP-element group 46: 	 branch_block_stmt_655/if_stmt_832_if_link/if_choice_transition
      -- CP-element group 46: 	 branch_block_stmt_655/lorx_xlhsx_xfalse48_ifx_xthen
      -- CP-element group 46: 	 branch_block_stmt_655/lorx_xlhsx_xfalse48_ifx_xthen_PhiReq/$entry
      -- CP-element group 46: 	 branch_block_stmt_655/lorx_xlhsx_xfalse48_ifx_xthen_PhiReq/$exit
      -- 
    if_choice_transition_2916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_832_branch_ack_1, ack => zeropad3D_CP_2067_elements(46)); -- 
    -- CP-element group 47:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	49 
    -- CP-element group 47: 	51 
    -- CP-element group 47:  members (27) 
      -- CP-element group 47: 	 branch_block_stmt_655/merge_stmt_838__exit__
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863__entry__
      -- CP-element group 47: 	 branch_block_stmt_655/if_stmt_832_else_link/$exit
      -- CP-element group 47: 	 branch_block_stmt_655/if_stmt_832_else_link/else_choice_transition
      -- CP-element group 47: 	 branch_block_stmt_655/lorx_xlhsx_xfalse48_lorx_xlhsx_xfalse55
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_update_start_
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_word_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Sample/word_access_start/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Sample/word_access_start/word_0/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Sample/word_access_start/word_0/rr
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/word_access_complete/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/word_access_complete/word_0/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/word_access_complete/word_0/cr
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_update_start_
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_Update/cr
      -- CP-element group 47: 	 branch_block_stmt_655/lorx_xlhsx_xfalse48_lorx_xlhsx_xfalse55_PhiReq/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/lorx_xlhsx_xfalse48_lorx_xlhsx_xfalse55_PhiReq/$exit
      -- CP-element group 47: 	 branch_block_stmt_655/merge_stmt_838_PhiReqMerge
      -- CP-element group 47: 	 branch_block_stmt_655/merge_stmt_838_PhiAck/$entry
      -- CP-element group 47: 	 branch_block_stmt_655/merge_stmt_838_PhiAck/$exit
      -- CP-element group 47: 	 branch_block_stmt_655/merge_stmt_838_PhiAck/dummy
      -- 
    else_choice_transition_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_832_branch_ack_0, ack => zeropad3D_CP_2067_elements(47)); -- 
    rr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(47), ack => LOAD_col_high_840_load_0_req_0); -- 
    cr_2952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(47), ack => LOAD_col_high_840_load_0_req_1); -- 
    cr_2971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(47), ack => type_cast_844_inst_req_1); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Sample/word_access_start/$exit
      -- CP-element group 48: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Sample/word_access_start/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Sample/word_access_start/word_0/ra
      -- 
    ra_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_840_load_0_ack_0, ack => zeropad3D_CP_2067_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (12) 
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/word_access_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/word_access_complete/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/word_access_complete/word_0/ca
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/LOAD_col_high_840_Merge/$entry
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/LOAD_col_high_840_Merge/$exit
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/LOAD_col_high_840_Merge/merge_req
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/LOAD_col_high_840_Update/LOAD_col_high_840_Merge/merge_ack
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_Sample/rr
      -- 
    ca_2953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_840_load_0_ack_1, ack => zeropad3D_CP_2067_elements(49)); -- 
    rr_2966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(49), ack => type_cast_844_inst_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_Sample/ra
      -- 
    ra_2967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_844_inst_ack_0, ack => zeropad3D_CP_2067_elements(50)); -- 
    -- CP-element group 51:  branch  transition  place  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	47 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863__exit__
      -- CP-element group 51: 	 branch_block_stmt_655/if_stmt_864__entry__
      -- CP-element group 51: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/$exit
      -- CP-element group 51: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_655/assign_stmt_841_to_assign_stmt_863/type_cast_844_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_655/if_stmt_864_dead_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_655/if_stmt_864_eval_test/$entry
      -- CP-element group 51: 	 branch_block_stmt_655/if_stmt_864_eval_test/$exit
      -- CP-element group 51: 	 branch_block_stmt_655/if_stmt_864_eval_test/branch_req
      -- CP-element group 51: 	 branch_block_stmt_655/R_cmp64_865_place
      -- CP-element group 51: 	 branch_block_stmt_655/if_stmt_864_if_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_655/if_stmt_864_else_link/$entry
      -- 
    ca_2972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_844_inst_ack_1, ack => zeropad3D_CP_2067_elements(51)); -- 
    branch_req_2980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(51), ack => if_stmt_864_branch_req_0); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52: 	69 
    -- CP-element group 52: 	71 
    -- CP-element group 52: 	73 
    -- CP-element group 52: 	75 
    -- CP-element group 52: 	77 
    -- CP-element group 52: 	79 
    -- CP-element group 52: 	81 
    -- CP-element group 52: 	83 
    -- CP-element group 52: 	86 
    -- CP-element group 52:  members (46) 
      -- CP-element group 52: 	 branch_block_stmt_655/merge_stmt_929__exit__
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034__entry__
      -- CP-element group 52: 	 branch_block_stmt_655/if_stmt_864_if_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_655/if_stmt_864_if_link/if_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_655/lorx_xlhsx_xfalse55_ifx_xelse
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_update_start_
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_update_start_
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_update_start_
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_update_start
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_Update/req
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_complete/req
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_update_start_
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_update_start_
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_update_start_
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_update_start
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_Update/req
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_complete/req
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_update_start_
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_655/lorx_xlhsx_xfalse55_ifx_xelse_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/lorx_xlhsx_xfalse55_ifx_xelse_PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_655/merge_stmt_929_PhiReqMerge
      -- CP-element group 52: 	 branch_block_stmt_655/merge_stmt_929_PhiAck/$entry
      -- CP-element group 52: 	 branch_block_stmt_655/merge_stmt_929_PhiAck/$exit
      -- CP-element group 52: 	 branch_block_stmt_655/merge_stmt_929_PhiAck/dummy
      -- 
    if_choice_transition_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_864_branch_ack_1, ack => zeropad3D_CP_2067_elements(52)); -- 
    rr_3143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => type_cast_933_inst_req_0); -- 
    cr_3148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => type_cast_933_inst_req_1); -- 
    cr_3162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => type_cast_997_inst_req_1); -- 
    req_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => array_obj_ref_1003_index_offset_req_1); -- 
    req_3208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => addr_of_1004_final_reg_req_1); -- 
    cr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => ptr_deref_1008_load_0_req_1); -- 
    cr_3272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => type_cast_1022_inst_req_1); -- 
    req_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => array_obj_ref_1028_index_offset_req_1); -- 
    req_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => addr_of_1029_final_reg_req_1); -- 
    cr_3368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(52), ack => ptr_deref_1032_store_0_req_1); -- 
    -- CP-element group 53:  transition  place  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	816 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_655/if_stmt_864_else_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_655/if_stmt_864_else_link/else_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_655/lorx_xlhsx_xfalse55_ifx_xthen
      -- CP-element group 53: 	 branch_block_stmt_655/lorx_xlhsx_xfalse55_ifx_xthen_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_655/lorx_xlhsx_xfalse55_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_864_branch_ack_0, ack => zeropad3D_CP_2067_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	816 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_Sample/ra
      -- 
    ra_3003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_874_inst_ack_0, ack => zeropad3D_CP_2067_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	816 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_Update/ca
      -- 
    ca_3008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_874_inst_ack_1, ack => zeropad3D_CP_2067_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	816 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_Sample/ra
      -- 
    ra_3017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_879_inst_ack_0, ack => zeropad3D_CP_2067_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	816 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_Update/ca
      -- 
    ca_3022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_879_inst_ack_1, ack => zeropad3D_CP_2067_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_Sample/rr
      -- 
    rr_3030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(58), ack => type_cast_914_inst_req_0); -- 
    zeropad3D_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(57) & zeropad3D_CP_2067_elements(55);
      gj_zeropad3D_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_Sample/ra
      -- 
    ra_3031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_914_inst_ack_0, ack => zeropad3D_CP_2067_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	816 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (16) 
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_resized_1
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_scaled_1
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_computed_1
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_resize_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_resize_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_resize_1/index_resize_req
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_resize_1/index_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_scale_1/$entry
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_scale_1/$exit
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_scale_1/scale_rename_req
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_index_scale_1/scale_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_Sample/req
      -- 
    ca_3036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_914_inst_ack_1, ack => zeropad3D_CP_2067_elements(60)); -- 
    req_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(60), ack => array_obj_ref_920_index_offset_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	67 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_sample_complete
      -- CP-element group 61: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_Sample/ack
      -- 
    ack_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_920_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	816 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (11) 
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_offset_calculated
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_request/$entry
      -- CP-element group 62: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_request/req
      -- 
    ack_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_920_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(62)); -- 
    req_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(62), ack => addr_of_921_final_reg_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_request/$exit
      -- CP-element group 63: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_request/ack
      -- 
    ack_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_921_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	816 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (28) 
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_complete/ack
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_word_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_root_address_calculated
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_address_resized
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_addr_resize/$entry
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_addr_resize/$exit
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_addr_resize/base_resize_req
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_addr_resize/base_resize_ack
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_plus_offset/$entry
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_plus_offset/$exit
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_plus_offset/sum_rename_req
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_base_plus_offset/sum_rename_ack
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_word_addrgen/$entry
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_word_addrgen/$exit
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_word_addrgen/root_register_req
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_word_addrgen/root_register_ack
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/ptr_deref_924_Split/$entry
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/ptr_deref_924_Split/$exit
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/ptr_deref_924_Split/split_req
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/ptr_deref_924_Split/split_ack
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/word_access_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/word_access_start/word_0/$entry
      -- CP-element group 64: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/word_access_start/word_0/rr
      -- 
    ack_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_921_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(64)); -- 
    rr_3120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(64), ack => ptr_deref_924_store_0_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/word_access_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/word_access_start/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Sample/word_access_start/word_0/ra
      -- 
    ra_3121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_924_store_0_ack_0, ack => zeropad3D_CP_2067_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	816 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Update/word_access_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Update/word_access_complete/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Update/word_access_complete/word_0/ca
      -- 
    ca_3132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_924_store_0_ack_1, ack => zeropad3D_CP_2067_elements(66)); -- 
    -- CP-element group 67:  join  transition  place  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	61 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	817 
    -- CP-element group 67:  members (5) 
      -- CP-element group 67: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927__exit__
      -- CP-element group 67: 	 branch_block_stmt_655/ifx_xthen_ifx_xend
      -- CP-element group 67: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/$exit
      -- CP-element group 67: 	 branch_block_stmt_655/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_655/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(61) & zeropad3D_CP_2067_elements(66);
      gj_zeropad3D_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_Sample/ra
      -- 
    ra_3144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_933_inst_ack_0, ack => zeropad3D_CP_2067_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	52 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: 	78 
    -- CP-element group 69:  members (9) 
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_933_Update/ca
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_Sample/rr
      -- 
    ca_3149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_933_inst_ack_1, ack => zeropad3D_CP_2067_elements(69)); -- 
    rr_3157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(69), ack => type_cast_997_inst_req_0); -- 
    rr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(69), ack => type_cast_1022_inst_req_0); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_Sample/ra
      -- 
    ra_3158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_997_inst_ack_0, ack => zeropad3D_CP_2067_elements(70)); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	52 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (16) 
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_997_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_resized_1
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_scaled_1
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_computed_1
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_resize_1/$entry
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_resize_1/$exit
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_resize_1/index_resize_req
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_resize_1/index_resize_ack
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_scale_1/$entry
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_scale_1/$exit
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_scale_1/scale_rename_req
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_index_scale_1/scale_rename_ack
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_Sample/req
      -- 
    ca_3163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_997_inst_ack_1, ack => zeropad3D_CP_2067_elements(71)); -- 
    req_3188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(71), ack => array_obj_ref_1003_index_offset_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	87 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_sample_complete
      -- CP-element group 72: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_Sample/ack
      -- 
    ack_3189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1003_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(72)); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	52 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (11) 
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_offset_calculated
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_final_index_sum_regn_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1003_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_request/$entry
      -- CP-element group 73: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_request/req
      -- 
    ack_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1003_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(73)); -- 
    req_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(73), ack => addr_of_1004_final_reg_req_0); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_request/$exit
      -- CP-element group 74: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_request/ack
      -- 
    ack_3204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1004_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (24) 
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1004_complete/ack
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_word_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_root_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_address_resized
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_addr_resize/$entry
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_addr_resize/$exit
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_addr_resize/base_resize_req
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_addr_resize/base_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_plus_offset/$entry
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_plus_offset/$exit
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_plus_offset/sum_rename_req
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_base_plus_offset/sum_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_word_addrgen/$entry
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_word_addrgen/$exit
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_word_addrgen/root_register_req
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_word_addrgen/root_register_ack
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Sample/word_access_start/$entry
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Sample/word_access_start/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Sample/word_access_start/word_0/rr
      -- 
    ack_3209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1004_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(75)); -- 
    rr_3242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(75), ack => ptr_deref_1008_load_0_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Sample/word_access_start/$exit
      -- CP-element group 76: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Sample/word_access_start/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Sample/word_access_start/word_0/ra
      -- 
    ra_3243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1008_load_0_ack_0, ack => zeropad3D_CP_2067_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	52 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	84 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/word_access_complete/$exit
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/word_access_complete/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/word_access_complete/word_0/ca
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/ptr_deref_1008_Merge/$entry
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/ptr_deref_1008_Merge/$exit
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/ptr_deref_1008_Merge/merge_req
      -- CP-element group 77: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1008_Update/ptr_deref_1008_Merge/merge_ack
      -- 
    ca_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1008_load_0_ack_1, ack => zeropad3D_CP_2067_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	69 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_Sample/ra
      -- 
    ra_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1022_inst_ack_0, ack => zeropad3D_CP_2067_elements(78)); -- 
    -- CP-element group 79:  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	52 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (16) 
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/type_cast_1022_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_resized_1
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_scaled_1
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_computed_1
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_resize_1/$entry
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_resize_1/$exit
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_resize_1/index_resize_req
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_resize_1/index_resize_ack
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_scale_1/$entry
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_scale_1/$exit
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_scale_1/scale_rename_req
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_index_scale_1/scale_rename_ack
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_Sample/req
      -- 
    ca_3273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1022_inst_ack_1, ack => zeropad3D_CP_2067_elements(79)); -- 
    req_3298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(79), ack => array_obj_ref_1028_index_offset_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	87 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_sample_complete
      -- CP-element group 80: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_Sample/ack
      -- 
    ack_3299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	52 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (11) 
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_root_address_calculated
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_offset_calculated
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_final_index_sum_regn_Update/ack
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_base_plus_offset/$entry
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_base_plus_offset/$exit
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_base_plus_offset/sum_rename_req
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/array_obj_ref_1028_base_plus_offset/sum_rename_ack
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_request/$entry
      -- CP-element group 81: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_request/req
      -- 
    ack_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(81)); -- 
    req_3313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(81), ack => addr_of_1029_final_reg_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_request/$exit
      -- CP-element group 82: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_request/ack
      -- 
    ack_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1029_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	52 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (19) 
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_complete/$exit
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/addr_of_1029_complete/ack
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_address_calculated
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_word_address_calculated
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_root_address_calculated
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_address_resized
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_addr_resize/$entry
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_addr_resize/$exit
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_addr_resize/base_resize_req
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_addr_resize/base_resize_ack
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_plus_offset/$entry
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_plus_offset/$exit
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_plus_offset/sum_rename_req
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_base_plus_offset/sum_rename_ack
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_word_addrgen/$entry
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_word_addrgen/$exit
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_word_addrgen/root_register_req
      -- CP-element group 83: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_word_addrgen/root_register_ack
      -- 
    ack_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1029_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	77 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/ptr_deref_1032_Split/$entry
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/ptr_deref_1032_Split/$exit
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/ptr_deref_1032_Split/split_req
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/ptr_deref_1032_Split/split_ack
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/word_access_start/$entry
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/word_access_start/word_0/$entry
      -- CP-element group 84: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/word_access_start/word_0/rr
      -- 
    rr_3357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(84), ack => ptr_deref_1032_store_0_req_0); -- 
    zeropad3D_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(77) & zeropad3D_CP_2067_elements(83);
      gj_zeropad3D_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/word_access_start/$exit
      -- CP-element group 85: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/word_access_start/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Sample/word_access_start/word_0/ra
      -- 
    ra_3358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1032_store_0_ack_0, ack => zeropad3D_CP_2067_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	52 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Update/word_access_complete/$exit
      -- CP-element group 86: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Update/word_access_complete/word_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/ptr_deref_1032_Update/word_access_complete/word_0/ca
      -- 
    ca_3369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1032_store_0_ack_1, ack => zeropad3D_CP_2067_elements(86)); -- 
    -- CP-element group 87:  join  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	72 
    -- CP-element group 87: 	80 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	817 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034__exit__
      -- CP-element group 87: 	 branch_block_stmt_655/ifx_xelse_ifx_xend
      -- CP-element group 87: 	 branch_block_stmt_655/assign_stmt_934_to_assign_stmt_1034/$exit
      -- CP-element group 87: 	 branch_block_stmt_655/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_655/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(72) & zeropad3D_CP_2067_elements(80) & zeropad3D_CP_2067_elements(86);
      gj_zeropad3D_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	817 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_Sample/ra
      -- 
    ra_3381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1040_inst_ack_0, ack => zeropad3D_CP_2067_elements(88)); -- 
    -- CP-element group 89:  branch  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	817 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (13) 
      -- CP-element group 89: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054__exit__
      -- CP-element group 89: 	 branch_block_stmt_655/if_stmt_1055__entry__
      -- CP-element group 89: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/$exit
      -- CP-element group 89: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_655/if_stmt_1055_dead_link/$entry
      -- CP-element group 89: 	 branch_block_stmt_655/if_stmt_1055_eval_test/$entry
      -- CP-element group 89: 	 branch_block_stmt_655/if_stmt_1055_eval_test/$exit
      -- CP-element group 89: 	 branch_block_stmt_655/if_stmt_1055_eval_test/branch_req
      -- CP-element group 89: 	 branch_block_stmt_655/R_cmp133_1056_place
      -- CP-element group 89: 	 branch_block_stmt_655/if_stmt_1055_if_link/$entry
      -- CP-element group 89: 	 branch_block_stmt_655/if_stmt_1055_else_link/$entry
      -- 
    ca_3386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1040_inst_ack_1, ack => zeropad3D_CP_2067_elements(89)); -- 
    branch_req_3394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(89), ack => if_stmt_1055_branch_req_0); -- 
    -- CP-element group 90:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	826 
    -- CP-element group 90: 	827 
    -- CP-element group 90: 	829 
    -- CP-element group 90: 	830 
    -- CP-element group 90: 	832 
    -- CP-element group 90: 	833 
    -- CP-element group 90:  members (40) 
      -- CP-element group 90: 	 branch_block_stmt_655/merge_stmt_1061__exit__
      -- CP-element group 90: 	 branch_block_stmt_655/assign_stmt_1067__entry__
      -- CP-element group 90: 	 branch_block_stmt_655/assign_stmt_1067__exit__
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174
      -- CP-element group 90: 	 branch_block_stmt_655/if_stmt_1055_if_link/$exit
      -- CP-element group 90: 	 branch_block_stmt_655/if_stmt_1055_if_link/if_choice_transition
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xend_ifx_xthen135
      -- CP-element group 90: 	 branch_block_stmt_655/assign_stmt_1067/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/assign_stmt_1067/$exit
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xend_ifx_xthen135_PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xend_ifx_xthen135_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_655/merge_stmt_1061_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_655/merge_stmt_1061_PhiAck/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/merge_stmt_1061_PhiAck/$exit
      -- CP-element group 90: 	 branch_block_stmt_655/merge_stmt_1061_PhiAck/dummy
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/Update/cr
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Update/cr
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1055_branch_ack_1, ack => zeropad3D_CP_2067_elements(90)); -- 
    rr_10935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(90), ack => type_cast_1158_inst_req_0); -- 
    cr_10940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(90), ack => type_cast_1158_inst_req_1); -- 
    rr_10958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(90), ack => type_cast_1164_inst_req_0); -- 
    cr_10963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(90), ack => type_cast_1164_inst_req_1); -- 
    rr_10981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(90), ack => type_cast_1170_inst_req_0); -- 
    cr_10986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(90), ack => type_cast_1170_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  place  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	93 
    -- CP-element group 91: 	94 
    -- CP-element group 91: 	95 
    -- CP-element group 91: 	97 
    -- CP-element group 91: 	100 
    -- CP-element group 91: 	102 
    -- CP-element group 91: 	103 
    -- CP-element group 91: 	104 
    -- CP-element group 91: 	106 
    -- CP-element group 91:  members (54) 
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_update_start_
      -- CP-element group 91: 	 branch_block_stmt_655/merge_stmt_1069__exit__
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147__entry__
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/word_access_complete/word_0/cr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/word_access_complete/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/word_access_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Sample/word_access_start/word_0/rr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Sample/word_access_start/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Sample/word_access_start/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/if_stmt_1055_else_link/$exit
      -- CP-element group 91: 	 branch_block_stmt_655/if_stmt_1055_else_link/else_choice_transition
      -- CP-element group 91: 	 branch_block_stmt_655/ifx_xend_ifx_xelse140
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_update_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_update_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_word_address_calculated
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_root_address_calculated
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Sample/word_access_start/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Sample/word_access_start/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Sample/word_access_start/word_0/rr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/word_access_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/word_access_complete/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/word_access_complete/word_0/cr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_update_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_update_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_update_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_update_start_
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_word_address_calculated
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_root_address_calculated
      -- CP-element group 91: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/ifx_xend_ifx_xelse140_PhiReq/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/ifx_xend_ifx_xelse140_PhiReq/$exit
      -- CP-element group 91: 	 branch_block_stmt_655/merge_stmt_1069_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_655/merge_stmt_1069_PhiAck/$entry
      -- CP-element group 91: 	 branch_block_stmt_655/merge_stmt_1069_PhiAck/$exit
      -- CP-element group 91: 	 branch_block_stmt_655/merge_stmt_1069_PhiAck/dummy
      -- 
    else_choice_transition_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1055_branch_ack_0, ack => zeropad3D_CP_2067_elements(91)); -- 
    cr_3527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => LOAD_row_high_1126_load_0_req_1); -- 
    rr_3516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => LOAD_row_high_1126_load_0_req_0); -- 
    cr_3546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => type_cast_1130_inst_req_1); -- 
    rr_3419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => type_cast_1079_inst_req_0); -- 
    cr_3424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => type_cast_1079_inst_req_1); -- 
    rr_3441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => LOAD_col_high_1082_load_0_req_0); -- 
    cr_3452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => LOAD_col_high_1082_load_0_req_1); -- 
    cr_3471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => type_cast_1086_inst_req_1); -- 
    cr_3485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => type_cast_1106_inst_req_1); -- 
    cr_3499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(91), ack => type_cast_1123_inst_req_1); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_Sample/ra
      -- 
    ra_3420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1079_inst_ack_0, ack => zeropad3D_CP_2067_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	98 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1079_Update/ca
      -- 
    ca_3425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1079_inst_ack_1, ack => zeropad3D_CP_2067_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Sample/word_access_start/$exit
      -- CP-element group 94: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Sample/word_access_start/word_0/$exit
      -- CP-element group 94: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Sample/word_access_start/word_0/ra
      -- 
    ra_3442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1082_load_0_ack_0, ack => zeropad3D_CP_2067_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	91 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (12) 
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/word_access_complete/$exit
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/word_access_complete/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/word_access_complete/word_0/ca
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/LOAD_col_high_1082_Merge/$entry
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/LOAD_col_high_1082_Merge/$exit
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/LOAD_col_high_1082_Merge/merge_req
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_col_high_1082_Update/LOAD_col_high_1082_Merge/merge_ack
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_Sample/rr
      -- 
    ca_3453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1082_load_0_ack_1, ack => zeropad3D_CP_2067_elements(95)); -- 
    rr_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(95), ack => type_cast_1086_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_Sample/ra
      -- 
    ra_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1086_inst_ack_0, ack => zeropad3D_CP_2067_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	91 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1086_Update/ca
      -- 
    ca_3472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1086_inst_ack_1, ack => zeropad3D_CP_2067_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	93 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_Sample/rr
      -- 
    rr_3480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(98), ack => type_cast_1106_inst_req_0); -- 
    zeropad3D_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(93) & zeropad3D_CP_2067_elements(97);
      gj_zeropad3D_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_Sample/ra
      -- 
    ra_3481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_0, ack => zeropad3D_CP_2067_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	91 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1106_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_Sample/rr
      -- 
    ca_3486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_1, ack => zeropad3D_CP_2067_elements(100)); -- 
    rr_3494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(100), ack => type_cast_1123_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_Sample/ra
      -- 
    ra_3495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1123_inst_ack_0, ack => zeropad3D_CP_2067_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	91 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	107 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1123_Update/ca
      -- 
    ca_3500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1123_inst_ack_1, ack => zeropad3D_CP_2067_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	91 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Sample/word_access_start/word_0/ra
      -- CP-element group 103: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Sample/word_access_start/word_0/$exit
      -- CP-element group 103: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Sample/word_access_start/$exit
      -- CP-element group 103: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Sample/$exit
      -- 
    ra_3517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1126_load_0_ack_0, ack => zeropad3D_CP_2067_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	91 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (12) 
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/LOAD_row_high_1126_Merge/merge_ack
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/LOAD_row_high_1126_Merge/merge_req
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/LOAD_row_high_1126_Merge/$exit
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/LOAD_row_high_1126_Merge/$entry
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/word_access_complete/word_0/ca
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/word_access_complete/word_0/$exit
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/word_access_complete/$exit
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/LOAD_row_high_1126_update_completed_
      -- 
    ca_3528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1126_load_0_ack_1, ack => zeropad3D_CP_2067_elements(104)); -- 
    rr_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(104), ack => type_cast_1130_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_Sample/$exit
      -- 
    ra_3542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_0, ack => zeropad3D_CP_2067_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	91 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/type_cast_1130_Update/$exit
      -- 
    ca_3547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_1, ack => zeropad3D_CP_2067_elements(106)); -- 
    -- CP-element group 107:  branch  join  transition  place  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (10) 
      -- CP-element group 107: 	 branch_block_stmt_655/if_stmt_1148_else_link/$entry
      -- CP-element group 107: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147__exit__
      -- CP-element group 107: 	 branch_block_stmt_655/if_stmt_1148__entry__
      -- CP-element group 107: 	 branch_block_stmt_655/if_stmt_1148_if_link/$entry
      -- CP-element group 107: 	 branch_block_stmt_655/if_stmt_1148_eval_test/branch_req
      -- CP-element group 107: 	 branch_block_stmt_655/if_stmt_1148_eval_test/$exit
      -- CP-element group 107: 	 branch_block_stmt_655/if_stmt_1148_eval_test/$entry
      -- CP-element group 107: 	 branch_block_stmt_655/R_cmp166_1149_place
      -- CP-element group 107: 	 branch_block_stmt_655/if_stmt_1148_dead_link/$entry
      -- CP-element group 107: 	 branch_block_stmt_655/assign_stmt_1075_to_assign_stmt_1147/$exit
      -- 
    branch_req_3555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(107), ack => if_stmt_1148_branch_req_0); -- 
    zeropad3D_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(102) & zeropad3D_CP_2067_elements(106);
      gj_zeropad3D_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  fork  transition  place  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	841 
    -- CP-element group 108: 	842 
    -- CP-element group 108: 	844 
    -- CP-element group 108: 	845 
    -- CP-element group 108:  members (20) 
      -- CP-element group 108: 	 branch_block_stmt_655/if_stmt_1148_if_link/if_choice_transition
      -- CP-element group 108: 	 branch_block_stmt_655/if_stmt_1148_if_link/$exit
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/Update/cr
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1148_branch_ack_1, ack => zeropad3D_CP_2067_elements(108)); -- 
    rr_11014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(108), ack => type_cast_1180_inst_req_0); -- 
    cr_11019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(108), ack => type_cast_1180_inst_req_1); -- 
    rr_11037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(108), ack => type_cast_1184_inst_req_0); -- 
    cr_11042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(108), ack => type_cast_1184_inst_req_1); -- 
    -- CP-element group 109:  fork  transition  place  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	818 
    -- CP-element group 109: 	819 
    -- CP-element group 109: 	821 
    -- CP-element group 109: 	822 
    -- CP-element group 109: 	824 
    -- CP-element group 109:  members (22) 
      -- CP-element group 109: 	 branch_block_stmt_655/if_stmt_1148_else_link/$exit
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174
      -- CP-element group 109: 	 branch_block_stmt_655/if_stmt_1148_else_link/else_choice_transition
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/Update/cr
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/Update/cr
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1167/$entry
      -- CP-element group 109: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/$entry
      -- 
    else_choice_transition_3564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1148_branch_ack_0, ack => zeropad3D_CP_2067_elements(109)); -- 
    rr_10878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(109), ack => type_cast_1160_inst_req_0); -- 
    cr_10883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(109), ack => type_cast_1160_inst_req_1); -- 
    rr_10901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(109), ack => type_cast_1166_inst_req_0); -- 
    cr_10906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(109), ack => type_cast_1166_inst_req_1); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	850 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_Sample/ra
      -- 
    ra_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1188_inst_ack_0, ack => zeropad3D_CP_2067_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	850 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	130 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_Update/$exit
      -- 
    ca_3583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1188_inst_ack_1, ack => zeropad3D_CP_2067_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	850 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Sample/word_access_start/word_0/ra
      -- CP-element group 112: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Sample/word_access_start/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Sample/word_access_start/$exit
      -- CP-element group 112: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_sample_completed_
      -- 
    ra_3600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1197_load_0_ack_0, ack => zeropad3D_CP_2067_elements(112)); -- 
    -- CP-element group 113:  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	850 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	126 
    -- CP-element group 113:  members (12) 
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/LOAD_pad_1197_Merge/merge_ack
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/LOAD_pad_1197_Merge/merge_req
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/LOAD_pad_1197_Merge/$exit
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/LOAD_pad_1197_Merge/$entry
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/word_access_complete/word_0/ca
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/word_access_complete/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/word_access_complete/$exit
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_update_completed_
      -- 
    ca_3611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1197_load_0_ack_1, ack => zeropad3D_CP_2067_elements(113)); -- 
    rr_3765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(113), ack => type_cast_1227_inst_req_0); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	850 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Sample/word_access_start/word_0/ra
      -- CP-element group 114: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Sample/word_access_start/word_0/$exit
      -- CP-element group 114: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Sample/word_access_start/$exit
      -- CP-element group 114: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_sample_completed_
      -- 
    ra_3633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1200_load_0_ack_0, ack => zeropad3D_CP_2067_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	850 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	120 
    -- CP-element group 115:  members (12) 
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/LOAD_depth_high_1200_Merge/merge_ack
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/LOAD_depth_high_1200_Merge/merge_req
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/LOAD_depth_high_1200_Merge/$exit
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/LOAD_depth_high_1200_Merge/$entry
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/word_access_complete/word_0/ca
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/word_access_complete/word_0/$exit
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/word_access_complete/$exit
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_sample_start_
      -- 
    ca_3644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1200_load_0_ack_1, ack => zeropad3D_CP_2067_elements(115)); -- 
    rr_3723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(115), ack => type_cast_1210_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	850 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Sample/word_access_start/word_0/$exit
      -- CP-element group 116: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Sample/word_access_start/$exit
      -- CP-element group 116: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Sample/word_access_start/word_0/ra
      -- 
    ra_3666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_1203_load_0_ack_0, ack => zeropad3D_CP_2067_elements(116)); -- 
    -- CP-element group 117:  fork  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	850 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	122 
    -- CP-element group 117: 	128 
    -- CP-element group 117:  members (15) 
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/LOAD_out_depth_high_1203_Merge/merge_ack
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/LOAD_out_depth_high_1203_Merge/merge_req
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/LOAD_out_depth_high_1203_Merge/$exit
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/LOAD_out_depth_high_1203_Merge/$entry
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/word_access_complete/word_0/ca
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/word_access_complete/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/word_access_complete/$exit
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_sample_start_
      -- 
    ca_3677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_1203_load_0_ack_1, ack => zeropad3D_CP_2067_elements(117)); -- 
    rr_3737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(117), ack => type_cast_1214_inst_req_0); -- 
    rr_3779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(117), ack => type_cast_1231_inst_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	850 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Sample/word_access_start/word_0/ra
      -- CP-element group 118: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Sample/word_access_start/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Sample/word_access_start/$exit
      -- CP-element group 118: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Sample/$exit
      -- 
    ra_3699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_1206_load_0_ack_0, ack => zeropad3D_CP_2067_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	850 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (12) 
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/LOAD_out_col_high_1206_Merge/merge_ack
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/LOAD_out_col_high_1206_Merge/merge_req
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/LOAD_out_col_high_1206_Merge/$exit
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/LOAD_out_col_high_1206_Merge/$entry
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/word_access_complete/word_0/ca
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/word_access_complete/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/word_access_complete/$exit
      -- CP-element group 119: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/$exit
      -- 
    ca_3710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_1206_load_0_ack_1, ack => zeropad3D_CP_2067_elements(119)); -- 
    rr_3751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(119), ack => type_cast_1218_inst_req_0); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	115 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_sample_completed_
      -- 
    ra_3724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_0, ack => zeropad3D_CP_2067_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	850 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	130 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_Update/ca
      -- CP-element group 121: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_Update/$exit
      -- 
    ca_3729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_1, ack => zeropad3D_CP_2067_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	117 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_sample_completed_
      -- 
    ra_3738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1214_inst_ack_0, ack => zeropad3D_CP_2067_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	850 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	130 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_Update/$exit
      -- 
    ca_3743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1214_inst_ack_1, ack => zeropad3D_CP_2067_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_Sample/ra
      -- CP-element group 124: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_sample_completed_
      -- 
    ra_3752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_0, ack => zeropad3D_CP_2067_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	850 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	130 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_Update/$exit
      -- 
    ca_3757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_1, ack => zeropad3D_CP_2067_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	113 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_Sample/ra
      -- CP-element group 126: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_sample_completed_
      -- 
    ra_3766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1227_inst_ack_0, ack => zeropad3D_CP_2067_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	850 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	130 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_update_completed_
      -- 
    ca_3771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1227_inst_ack_1, ack => zeropad3D_CP_2067_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	117 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_Sample/ra
      -- CP-element group 128: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_sample_completed_
      -- 
    ra_3780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_0, ack => zeropad3D_CP_2067_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	850 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_Update/ca
      -- CP-element group 129: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_update_completed_
      -- 
    ca_3785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_1, ack => zeropad3D_CP_2067_elements(129)); -- 
    -- CP-element group 130:  join  fork  transition  place  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	111 
    -- CP-element group 130: 	121 
    -- CP-element group 130: 	123 
    -- CP-element group 130: 	125 
    -- CP-element group 130: 	127 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	861 
    -- CP-element group 130: 	862 
    -- CP-element group 130: 	864 
    -- CP-element group 130: 	865 
    -- CP-element group 130:  members (16) 
      -- CP-element group 130: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273__exit__
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234
      -- CP-element group 130: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/$exit
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/Update/cr
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1282/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1289/$entry
      -- CP-element group 130: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/$entry
      -- 
    rr_11141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(130), ack => type_cast_1279_inst_req_0); -- 
    cr_11146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(130), ack => type_cast_1279_inst_req_1); -- 
    zeropad3D_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(111) & zeropad3D_CP_2067_elements(121) & zeropad3D_CP_2067_elements(123) & zeropad3D_CP_2067_elements(125) & zeropad3D_CP_2067_elements(127) & zeropad3D_CP_2067_elements(129);
      gj_zeropad3D_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	871 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_sample_completed_
      -- 
    ra_3797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1300_inst_ack_0, ack => zeropad3D_CP_2067_elements(131)); -- 
    -- CP-element group 132:  branch  transition  place  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	871 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (13) 
      -- CP-element group 132: 	 branch_block_stmt_655/if_stmt_1309_eval_test/branch_req
      -- CP-element group 132: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308__exit__
      -- CP-element group 132: 	 branch_block_stmt_655/if_stmt_1309__entry__
      -- CP-element group 132: 	 branch_block_stmt_655/if_stmt_1309_eval_test/$exit
      -- CP-element group 132: 	 branch_block_stmt_655/if_stmt_1309_eval_test/$entry
      -- CP-element group 132: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_655/if_stmt_1309_dead_link/$entry
      -- CP-element group 132: 	 branch_block_stmt_655/if_stmt_1309_if_link/$entry
      -- CP-element group 132: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_655/R_cmp239_1310_place
      -- CP-element group 132: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/$exit
      -- CP-element group 132: 	 branch_block_stmt_655/if_stmt_1309_else_link/$entry
      -- 
    ca_3802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1300_inst_ack_1, ack => zeropad3D_CP_2067_elements(132)); -- 
    branch_req_3810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(132), ack => if_stmt_1309_branch_req_0); -- 
    -- CP-element group 133:  transition  place  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	872 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_655/if_stmt_1309_if_link/$exit
      -- CP-element group 133: 	 branch_block_stmt_655/whilex_xbody234_ifx_xthen269
      -- CP-element group 133: 	 branch_block_stmt_655/if_stmt_1309_if_link/if_choice_transition
      -- CP-element group 133: 	 branch_block_stmt_655/whilex_xbody234_ifx_xthen269_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_655/whilex_xbody234_ifx_xthen269_PhiReq/$exit
      -- 
    if_choice_transition_3815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1309_branch_ack_1, ack => zeropad3D_CP_2067_elements(133)); -- 
    -- CP-element group 134:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	136 
    -- CP-element group 134: 	138 
    -- CP-element group 134:  members (27) 
      -- CP-element group 134: 	 branch_block_stmt_655/merge_stmt_1315__exit__
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340__entry__
      -- CP-element group 134: 	 branch_block_stmt_655/whilex_xbody234_lorx_xlhsx_xfalse241
      -- CP-element group 134: 	 branch_block_stmt_655/if_stmt_1309_else_link/$exit
      -- CP-element group 134: 	 branch_block_stmt_655/if_stmt_1309_else_link/else_choice_transition
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_update_start_
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_word_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_root_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Sample/word_access_start/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Sample/word_access_start/word_0/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Sample/word_access_start/word_0/rr
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/word_access_complete/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/word_access_complete/word_0/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/word_access_complete/word_0/cr
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_update_start_
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_Update/cr
      -- CP-element group 134: 	 branch_block_stmt_655/whilex_xbody234_lorx_xlhsx_xfalse241_PhiReq/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/whilex_xbody234_lorx_xlhsx_xfalse241_PhiReq/$exit
      -- CP-element group 134: 	 branch_block_stmt_655/merge_stmt_1315_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_655/merge_stmt_1315_PhiAck/$entry
      -- CP-element group 134: 	 branch_block_stmt_655/merge_stmt_1315_PhiAck/$exit
      -- CP-element group 134: 	 branch_block_stmt_655/merge_stmt_1315_PhiAck/dummy
      -- 
    else_choice_transition_3819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1309_branch_ack_0, ack => zeropad3D_CP_2067_elements(134)); -- 
    rr_3840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(134), ack => LOAD_row_high_1317_load_0_req_0); -- 
    cr_3851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(134), ack => LOAD_row_high_1317_load_0_req_1); -- 
    cr_3870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(134), ack => type_cast_1321_inst_req_1); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Sample/word_access_start/$exit
      -- CP-element group 135: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Sample/word_access_start/word_0/$exit
      -- CP-element group 135: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Sample/word_access_start/word_0/ra
      -- 
    ra_3841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1317_load_0_ack_0, ack => zeropad3D_CP_2067_elements(135)); -- 
    -- CP-element group 136:  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (12) 
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/word_access_complete/$exit
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/word_access_complete/word_0/$exit
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/word_access_complete/word_0/ca
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/LOAD_row_high_1317_Merge/$entry
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/LOAD_row_high_1317_Merge/$exit
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/LOAD_row_high_1317_Merge/merge_req
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/LOAD_row_high_1317_Update/LOAD_row_high_1317_Merge/merge_ack
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_Sample/rr
      -- 
    ca_3852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1317_load_0_ack_1, ack => zeropad3D_CP_2067_elements(136)); -- 
    rr_3865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(136), ack => type_cast_1321_inst_req_0); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_Sample/ra
      -- 
    ra_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_0, ack => zeropad3D_CP_2067_elements(137)); -- 
    -- CP-element group 138:  branch  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	134 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (13) 
      -- CP-element group 138: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340__exit__
      -- CP-element group 138: 	 branch_block_stmt_655/if_stmt_1341__entry__
      -- CP-element group 138: 	 branch_block_stmt_655/R_cmp250_1342_place
      -- CP-element group 138: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/$exit
      -- CP-element group 138: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_655/assign_stmt_1318_to_assign_stmt_1340/type_cast_1321_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_655/if_stmt_1341_dead_link/$entry
      -- CP-element group 138: 	 branch_block_stmt_655/if_stmt_1341_eval_test/$entry
      -- CP-element group 138: 	 branch_block_stmt_655/if_stmt_1341_eval_test/$exit
      -- CP-element group 138: 	 branch_block_stmt_655/if_stmt_1341_eval_test/branch_req
      -- CP-element group 138: 	 branch_block_stmt_655/if_stmt_1341_if_link/$entry
      -- CP-element group 138: 	 branch_block_stmt_655/if_stmt_1341_else_link/$entry
      -- 
    ca_3871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_1, ack => zeropad3D_CP_2067_elements(138)); -- 
    branch_req_3879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(138), ack => if_stmt_1341_branch_req_0); -- 
    -- CP-element group 139:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: 	142 
    -- CP-element group 139:  members (18) 
      -- CP-element group 139: 	 branch_block_stmt_655/lorx_xlhsx_xfalse241_lorx_xlhsx_xfalse252
      -- CP-element group 139: 	 branch_block_stmt_655/merge_stmt_1347__exit__
      -- CP-element group 139: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359__entry__
      -- CP-element group 139: 	 branch_block_stmt_655/if_stmt_1341_if_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_655/if_stmt_1341_if_link/if_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/$entry
      -- CP-element group 139: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_update_start_
      -- CP-element group 139: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_Update/cr
      -- CP-element group 139: 	 branch_block_stmt_655/lorx_xlhsx_xfalse241_lorx_xlhsx_xfalse252_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_655/lorx_xlhsx_xfalse241_lorx_xlhsx_xfalse252_PhiReq/$exit
      -- CP-element group 139: 	 branch_block_stmt_655/merge_stmt_1347_PhiReqMerge
      -- CP-element group 139: 	 branch_block_stmt_655/merge_stmt_1347_PhiAck/$entry
      -- CP-element group 139: 	 branch_block_stmt_655/merge_stmt_1347_PhiAck/$exit
      -- CP-element group 139: 	 branch_block_stmt_655/merge_stmt_1347_PhiAck/dummy
      -- 
    if_choice_transition_3884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1341_branch_ack_1, ack => zeropad3D_CP_2067_elements(139)); -- 
    rr_3901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(139), ack => type_cast_1351_inst_req_0); -- 
    cr_3906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(139), ack => type_cast_1351_inst_req_1); -- 
    -- CP-element group 140:  transition  place  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	872 
    -- CP-element group 140:  members (5) 
      -- CP-element group 140: 	 branch_block_stmt_655/lorx_xlhsx_xfalse241_ifx_xthen269
      -- CP-element group 140: 	 branch_block_stmt_655/if_stmt_1341_else_link/$exit
      -- CP-element group 140: 	 branch_block_stmt_655/if_stmt_1341_else_link/else_choice_transition
      -- CP-element group 140: 	 branch_block_stmt_655/lorx_xlhsx_xfalse241_ifx_xthen269_PhiReq/$entry
      -- CP-element group 140: 	 branch_block_stmt_655/lorx_xlhsx_xfalse241_ifx_xthen269_PhiReq/$exit
      -- 
    else_choice_transition_3888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1341_branch_ack_0, ack => zeropad3D_CP_2067_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_Sample/ra
      -- 
    ra_3902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1351_inst_ack_0, ack => zeropad3D_CP_2067_elements(141)); -- 
    -- CP-element group 142:  branch  transition  place  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (13) 
      -- CP-element group 142: 	 branch_block_stmt_655/R_cmp257_1361_place
      -- CP-element group 142: 	 branch_block_stmt_655/if_stmt_1360_if_link/$entry
      -- CP-element group 142: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359__exit__
      -- CP-element group 142: 	 branch_block_stmt_655/if_stmt_1360__entry__
      -- CP-element group 142: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/$exit
      -- CP-element group 142: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_655/assign_stmt_1352_to_assign_stmt_1359/type_cast_1351_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_655/if_stmt_1360_dead_link/$entry
      -- CP-element group 142: 	 branch_block_stmt_655/if_stmt_1360_eval_test/$entry
      -- CP-element group 142: 	 branch_block_stmt_655/if_stmt_1360_eval_test/$exit
      -- CP-element group 142: 	 branch_block_stmt_655/if_stmt_1360_eval_test/branch_req
      -- CP-element group 142: 	 branch_block_stmt_655/if_stmt_1360_else_link/$entry
      -- 
    ca_3907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1351_inst_ack_1, ack => zeropad3D_CP_2067_elements(142)); -- 
    branch_req_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(142), ack => if_stmt_1360_branch_req_0); -- 
    -- CP-element group 143:  transition  place  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	872 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_655/if_stmt_1360_if_link/$exit
      -- CP-element group 143: 	 branch_block_stmt_655/if_stmt_1360_if_link/if_choice_transition
      -- CP-element group 143: 	 branch_block_stmt_655/lorx_xlhsx_xfalse252_ifx_xthen269
      -- CP-element group 143: 	 branch_block_stmt_655/lorx_xlhsx_xfalse252_ifx_xthen269_PhiReq/$entry
      -- CP-element group 143: 	 branch_block_stmt_655/lorx_xlhsx_xfalse252_ifx_xthen269_PhiReq/$exit
      -- 
    if_choice_transition_3920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1360_branch_ack_1, ack => zeropad3D_CP_2067_elements(143)); -- 
    -- CP-element group 144:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144: 	146 
    -- CP-element group 144: 	148 
    -- CP-element group 144:  members (27) 
      -- CP-element group 144: 	 branch_block_stmt_655/merge_stmt_1366__exit__
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385__entry__
      -- CP-element group 144: 	 branch_block_stmt_655/lorx_xlhsx_xfalse252_lorx_xlhsx_xfalse259
      -- CP-element group 144: 	 branch_block_stmt_655/if_stmt_1360_else_link/$exit
      -- CP-element group 144: 	 branch_block_stmt_655/if_stmt_1360_else_link/else_choice_transition
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_update_start_
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_word_address_calculated
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_root_address_calculated
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Sample/word_access_start/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Sample/word_access_start/word_0/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Sample/word_access_start/word_0/rr
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/word_access_complete/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/word_access_complete/word_0/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/word_access_complete/word_0/cr
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_update_start_
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_Update/cr
      -- CP-element group 144: 	 branch_block_stmt_655/lorx_xlhsx_xfalse252_lorx_xlhsx_xfalse259_PhiReq/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/lorx_xlhsx_xfalse252_lorx_xlhsx_xfalse259_PhiReq/$exit
      -- CP-element group 144: 	 branch_block_stmt_655/merge_stmt_1366_PhiReqMerge
      -- CP-element group 144: 	 branch_block_stmt_655/merge_stmt_1366_PhiAck/$entry
      -- CP-element group 144: 	 branch_block_stmt_655/merge_stmt_1366_PhiAck/$exit
      -- CP-element group 144: 	 branch_block_stmt_655/merge_stmt_1366_PhiAck/dummy
      -- 
    else_choice_transition_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1360_branch_ack_0, ack => zeropad3D_CP_2067_elements(144)); -- 
    rr_3945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(144), ack => LOAD_col_high_1368_load_0_req_0); -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(144), ack => LOAD_col_high_1368_load_0_req_1); -- 
    cr_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(144), ack => type_cast_1372_inst_req_1); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Sample/word_access_start/$exit
      -- CP-element group 145: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Sample/word_access_start/word_0/ra
      -- 
    ra_3946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1368_load_0_ack_0, ack => zeropad3D_CP_2067_elements(145)); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (12) 
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/word_access_complete/$exit
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/word_access_complete/word_0/$exit
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/word_access_complete/word_0/ca
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/LOAD_col_high_1368_Merge/$entry
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/LOAD_col_high_1368_Merge/$exit
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/LOAD_col_high_1368_Merge/merge_req
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/LOAD_col_high_1368_Update/LOAD_col_high_1368_Merge/merge_ack
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_Sample/rr
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1368_load_0_ack_1, ack => zeropad3D_CP_2067_elements(146)); -- 
    rr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(146), ack => type_cast_1372_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_Sample/ra
      -- 
    ra_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1372_inst_ack_0, ack => zeropad3D_CP_2067_elements(147)); -- 
    -- CP-element group 148:  branch  transition  place  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	144 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (13) 
      -- CP-element group 148: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385__exit__
      -- CP-element group 148: 	 branch_block_stmt_655/if_stmt_1386__entry__
      -- CP-element group 148: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/$exit
      -- CP-element group 148: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_655/assign_stmt_1369_to_assign_stmt_1385/type_cast_1372_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_655/if_stmt_1386_dead_link/$entry
      -- CP-element group 148: 	 branch_block_stmt_655/if_stmt_1386_eval_test/$entry
      -- CP-element group 148: 	 branch_block_stmt_655/if_stmt_1386_eval_test/$exit
      -- CP-element group 148: 	 branch_block_stmt_655/if_stmt_1386_eval_test/branch_req
      -- CP-element group 148: 	 branch_block_stmt_655/R_cmp267_1387_place
      -- CP-element group 148: 	 branch_block_stmt_655/if_stmt_1386_if_link/$entry
      -- CP-element group 148: 	 branch_block_stmt_655/if_stmt_1386_else_link/$entry
      -- 
    ca_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1372_inst_ack_1, ack => zeropad3D_CP_2067_elements(148)); -- 
    branch_req_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(148), ack => if_stmt_1386_branch_req_0); -- 
    -- CP-element group 149:  fork  transition  place  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	165 
    -- CP-element group 149: 	166 
    -- CP-element group 149: 	168 
    -- CP-element group 149: 	170 
    -- CP-element group 149: 	172 
    -- CP-element group 149: 	174 
    -- CP-element group 149: 	176 
    -- CP-element group 149: 	178 
    -- CP-element group 149: 	180 
    -- CP-element group 149: 	183 
    -- CP-element group 149:  members (46) 
      -- CP-element group 149: 	 branch_block_stmt_655/merge_stmt_1450__exit__
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555__entry__
      -- CP-element group 149: 	 branch_block_stmt_655/if_stmt_1386_if_link/$exit
      -- CP-element group 149: 	 branch_block_stmt_655/if_stmt_1386_if_link/if_choice_transition
      -- CP-element group 149: 	 branch_block_stmt_655/lorx_xlhsx_xfalse259_ifx_xelse290
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_update_start_
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_update_start_
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_update_start_
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_update_start
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_Update/req
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_complete/req
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_update_start_
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/word_access_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/word_access_complete/word_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/word_access_complete/word_0/cr
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_update_start_
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_update_start_
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_update_start
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_Update/req
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_complete/req
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_update_start_
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Update/word_access_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Update/word_access_complete/word_0/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Update/word_access_complete/word_0/cr
      -- CP-element group 149: 	 branch_block_stmt_655/merge_stmt_1450_PhiAck/dummy
      -- CP-element group 149: 	 branch_block_stmt_655/lorx_xlhsx_xfalse259_ifx_xelse290_PhiReq/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/lorx_xlhsx_xfalse259_ifx_xelse290_PhiReq/$exit
      -- CP-element group 149: 	 branch_block_stmt_655/merge_stmt_1450_PhiReqMerge
      -- CP-element group 149: 	 branch_block_stmt_655/merge_stmt_1450_PhiAck/$entry
      -- CP-element group 149: 	 branch_block_stmt_655/merge_stmt_1450_PhiAck/$exit
      -- 
    if_choice_transition_3989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1386_branch_ack_1, ack => zeropad3D_CP_2067_elements(149)); -- 
    rr_4147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => type_cast_1454_inst_req_0); -- 
    cr_4152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => type_cast_1454_inst_req_1); -- 
    cr_4166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => type_cast_1518_inst_req_1); -- 
    req_4197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => array_obj_ref_1524_index_offset_req_1); -- 
    req_4212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => addr_of_1525_final_reg_req_1); -- 
    cr_4257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => ptr_deref_1529_load_0_req_1); -- 
    cr_4276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => type_cast_1543_inst_req_1); -- 
    req_4307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => array_obj_ref_1549_index_offset_req_1); -- 
    req_4322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => addr_of_1550_final_reg_req_1); -- 
    cr_4372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(149), ack => ptr_deref_1553_store_0_req_1); -- 
    -- CP-element group 150:  transition  place  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	872 
    -- CP-element group 150:  members (5) 
      -- CP-element group 150: 	 branch_block_stmt_655/if_stmt_1386_else_link/$exit
      -- CP-element group 150: 	 branch_block_stmt_655/if_stmt_1386_else_link/else_choice_transition
      -- CP-element group 150: 	 branch_block_stmt_655/lorx_xlhsx_xfalse259_ifx_xthen269
      -- CP-element group 150: 	 branch_block_stmt_655/lorx_xlhsx_xfalse259_ifx_xthen269_PhiReq/$entry
      -- CP-element group 150: 	 branch_block_stmt_655/lorx_xlhsx_xfalse259_ifx_xthen269_PhiReq/$exit
      -- 
    else_choice_transition_3993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1386_branch_ack_0, ack => zeropad3D_CP_2067_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	872 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_Sample/ra
      -- 
    ra_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_0, ack => zeropad3D_CP_2067_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	872 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_Update/ca
      -- 
    ca_4012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_1, ack => zeropad3D_CP_2067_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	872 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_Sample/ra
      -- 
    ra_4021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1401_inst_ack_0, ack => zeropad3D_CP_2067_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	872 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_Update/ca
      -- 
    ca_4026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1401_inst_ack_1, ack => zeropad3D_CP_2067_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	152 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_Sample/rr
      -- 
    rr_4034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(155), ack => type_cast_1435_inst_req_0); -- 
    zeropad3D_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(152) & zeropad3D_CP_2067_elements(154);
      gj_zeropad3D_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_Sample/ra
      -- 
    ra_4035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1435_inst_ack_0, ack => zeropad3D_CP_2067_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	872 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (16) 
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_resized_1
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_scaled_1
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_computed_1
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_resize_1/$entry
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_resize_1/$exit
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_resize_1/index_resize_req
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_resize_1/index_resize_ack
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_scale_1/$entry
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_scale_1/$exit
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_scale_1/scale_rename_req
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_index_scale_1/scale_rename_ack
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_Sample/req
      -- 
    ca_4040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1435_inst_ack_1, ack => zeropad3D_CP_2067_elements(157)); -- 
    req_4065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(157), ack => array_obj_ref_1441_index_offset_req_0); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	164 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_sample_complete
      -- CP-element group 158: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_Sample/ack
      -- 
    ack_4066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1441_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(158)); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	872 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (11) 
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_root_address_calculated
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_offset_calculated
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_Update/ack
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_base_plus_offset/$entry
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_base_plus_offset/$exit
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_base_plus_offset/sum_rename_req
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_base_plus_offset/sum_rename_ack
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_request/$entry
      -- CP-element group 159: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_request/req
      -- 
    ack_4071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1441_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(159)); -- 
    req_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(159), ack => addr_of_1442_final_reg_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_request/$exit
      -- CP-element group 160: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_request/ack
      -- 
    ack_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1442_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(160)); -- 
    -- CP-element group 161:  join  fork  transition  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	872 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (28) 
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_complete/$exit
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_complete/ack
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_word_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_root_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_address_resized
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_addr_resize/$entry
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_addr_resize/$exit
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_addr_resize/base_resize_req
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_addr_resize/base_resize_ack
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_plus_offset/$entry
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_plus_offset/$exit
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_plus_offset/sum_rename_req
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_base_plus_offset/sum_rename_ack
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_word_addrgen/$entry
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_word_addrgen/$exit
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_word_addrgen/root_register_req
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_word_addrgen/root_register_ack
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/ptr_deref_1445_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/ptr_deref_1445_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/ptr_deref_1445_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/ptr_deref_1445_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/word_access_start/word_0/rr
      -- 
    ack_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1442_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(161)); -- 
    rr_4124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(161), ack => ptr_deref_1445_store_0_req_0); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Sample/word_access_start/word_0/ra
      -- 
    ra_4125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1445_store_0_ack_0, ack => zeropad3D_CP_2067_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	872 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Update/word_access_complete/word_0/ca
      -- 
    ca_4136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1445_store_0_ack_1, ack => zeropad3D_CP_2067_elements(163)); -- 
    -- CP-element group 164:  join  transition  place  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	158 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	873 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448__exit__
      -- CP-element group 164: 	 branch_block_stmt_655/ifx_xthen269_ifx_xend338
      -- CP-element group 164: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/$exit
      -- CP-element group 164: 	 branch_block_stmt_655/ifx_xthen269_ifx_xend338_PhiReq/$exit
      -- CP-element group 164: 	 branch_block_stmt_655/ifx_xthen269_ifx_xend338_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(158) & zeropad3D_CP_2067_elements(163);
      gj_zeropad3D_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	149 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_Sample/ra
      -- 
    ra_4148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1454_inst_ack_0, ack => zeropad3D_CP_2067_elements(165)); -- 
    -- CP-element group 166:  fork  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	149 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166: 	175 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1454_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_Sample/rr
      -- 
    ca_4153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1454_inst_ack_1, ack => zeropad3D_CP_2067_elements(166)); -- 
    rr_4161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(166), ack => type_cast_1518_inst_req_0); -- 
    rr_4271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(166), ack => type_cast_1543_inst_req_0); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_Sample/ra
      -- 
    ra_4162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1518_inst_ack_0, ack => zeropad3D_CP_2067_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	149 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (16) 
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1518_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_resized_1
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_scaled_1
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_computed_1
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_resize_1/$entry
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_resize_1/$exit
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_resize_1/index_resize_req
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_resize_1/index_resize_ack
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_scale_1/$entry
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_scale_1/$exit
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_scale_1/scale_rename_req
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_index_scale_1/scale_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_Sample/req
      -- 
    ca_4167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1518_inst_ack_1, ack => zeropad3D_CP_2067_elements(168)); -- 
    req_4192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(168), ack => array_obj_ref_1524_index_offset_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	184 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_sample_complete
      -- CP-element group 169: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_Sample/ack
      -- 
    ack_4193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1524_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	149 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1524_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_request/req
      -- 
    ack_4198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1524_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(170)); -- 
    req_4207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(170), ack => addr_of_1525_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_request/ack
      -- 
    ack_4208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1525_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(171)); -- 
    -- CP-element group 172:  join  fork  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	149 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (24) 
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1525_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_word_addrgen/root_register_ack
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Sample/word_access_start/$entry
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Sample/word_access_start/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Sample/word_access_start/word_0/rr
      -- 
    ack_4213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1525_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(172)); -- 
    rr_4246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(172), ack => ptr_deref_1529_load_0_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (5) 
      -- CP-element group 173: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Sample/word_access_start/$exit
      -- CP-element group 173: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Sample/word_access_start/word_0/$exit
      -- CP-element group 173: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Sample/word_access_start/word_0/ra
      -- 
    ra_4247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_load_0_ack_0, ack => zeropad3D_CP_2067_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	149 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	181 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/word_access_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/word_access_complete/word_0/$exit
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/word_access_complete/word_0/ca
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/ptr_deref_1529_Merge/$entry
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/ptr_deref_1529_Merge/$exit
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/ptr_deref_1529_Merge/merge_req
      -- CP-element group 174: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1529_Update/ptr_deref_1529_Merge/merge_ack
      -- 
    ca_4258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_load_0_ack_1, ack => zeropad3D_CP_2067_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	166 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_Sample/ra
      -- 
    ra_4272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1543_inst_ack_0, ack => zeropad3D_CP_2067_elements(175)); -- 
    -- CP-element group 176:  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	149 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (16) 
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/type_cast_1543_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_resized_1
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_scaled_1
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_computed_1
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_resize_1/$entry
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_resize_1/$exit
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_resize_1/index_resize_req
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_resize_1/index_resize_ack
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_scale_1/$entry
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_scale_1/$exit
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_scale_1/scale_rename_req
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_index_scale_1/scale_rename_ack
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_Sample/req
      -- 
    ca_4277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1543_inst_ack_1, ack => zeropad3D_CP_2067_elements(176)); -- 
    req_4302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(176), ack => array_obj_ref_1549_index_offset_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	184 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_sample_complete
      -- CP-element group 177: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_Sample/ack
      -- 
    ack_4303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1549_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(177)); -- 
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	149 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (11) 
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_root_address_calculated
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_offset_calculated
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_final_index_sum_regn_Update/ack
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_base_plus_offset/$entry
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_base_plus_offset/$exit
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_base_plus_offset/sum_rename_req
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/array_obj_ref_1549_base_plus_offset/sum_rename_ack
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_request/$entry
      -- CP-element group 178: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_request/req
      -- 
    ack_4308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1549_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(178)); -- 
    req_4317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(178), ack => addr_of_1550_final_reg_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_request/$exit
      -- CP-element group 179: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_request/ack
      -- 
    ack_4318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1550_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(179)); -- 
    -- CP-element group 180:  fork  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	149 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (19) 
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_complete/$exit
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/addr_of_1550_complete/ack
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_address_calculated
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_word_address_calculated
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_root_address_calculated
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_address_resized
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_addr_resize/$entry
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_addr_resize/$exit
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_addr_resize/base_resize_req
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_addr_resize/base_resize_ack
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_plus_offset/$entry
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_plus_offset/$exit
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_plus_offset/sum_rename_req
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_base_plus_offset/sum_rename_ack
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_word_addrgen/$entry
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_word_addrgen/$exit
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_word_addrgen/root_register_req
      -- CP-element group 180: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_word_addrgen/root_register_ack
      -- 
    ack_4323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1550_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	174 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (9) 
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/ptr_deref_1553_Split/$entry
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/ptr_deref_1553_Split/$exit
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/ptr_deref_1553_Split/split_req
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/ptr_deref_1553_Split/split_ack
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/word_access_start/$entry
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/word_access_start/word_0/$entry
      -- CP-element group 181: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/word_access_start/word_0/rr
      -- 
    rr_4361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(181), ack => ptr_deref_1553_store_0_req_0); -- 
    zeropad3D_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(174) & zeropad3D_CP_2067_elements(180);
      gj_zeropad3D_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/word_access_start/$exit
      -- CP-element group 182: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/word_access_start/word_0/$exit
      -- CP-element group 182: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Sample/word_access_start/word_0/ra
      -- 
    ra_4362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1553_store_0_ack_0, ack => zeropad3D_CP_2067_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	149 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (5) 
      -- CP-element group 183: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Update/word_access_complete/$exit
      -- CP-element group 183: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Update/word_access_complete/word_0/$exit
      -- CP-element group 183: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/ptr_deref_1553_Update/word_access_complete/word_0/ca
      -- 
    ca_4373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1553_store_0_ack_1, ack => zeropad3D_CP_2067_elements(183)); -- 
    -- CP-element group 184:  join  transition  place  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	169 
    -- CP-element group 184: 	177 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	873 
    -- CP-element group 184:  members (5) 
      -- CP-element group 184: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555__exit__
      -- CP-element group 184: 	 branch_block_stmt_655/ifx_xelse290_ifx_xend338
      -- CP-element group 184: 	 branch_block_stmt_655/assign_stmt_1455_to_assign_stmt_1555/$exit
      -- CP-element group 184: 	 branch_block_stmt_655/ifx_xelse290_ifx_xend338_PhiReq/$exit
      -- CP-element group 184: 	 branch_block_stmt_655/ifx_xelse290_ifx_xend338_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(169) & zeropad3D_CP_2067_elements(177) & zeropad3D_CP_2067_elements(183);
      gj_zeropad3D_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	873 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_Sample/ra
      -- 
    ra_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1561_inst_ack_0, ack => zeropad3D_CP_2067_elements(185)); -- 
    -- CP-element group 186:  branch  transition  place  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	873 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (13) 
      -- CP-element group 186: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575__exit__
      -- CP-element group 186: 	 branch_block_stmt_655/if_stmt_1576__entry__
      -- CP-element group 186: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/$exit
      -- CP-element group 186: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_655/if_stmt_1576_dead_link/$entry
      -- CP-element group 186: 	 branch_block_stmt_655/if_stmt_1576_eval_test/$entry
      -- CP-element group 186: 	 branch_block_stmt_655/if_stmt_1576_eval_test/$exit
      -- CP-element group 186: 	 branch_block_stmt_655/if_stmt_1576_eval_test/branch_req
      -- CP-element group 186: 	 branch_block_stmt_655/R_cmp346_1577_place
      -- CP-element group 186: 	 branch_block_stmt_655/if_stmt_1576_if_link/$entry
      -- CP-element group 186: 	 branch_block_stmt_655/if_stmt_1576_else_link/$entry
      -- 
    ca_4390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1561_inst_ack_1, ack => zeropad3D_CP_2067_elements(186)); -- 
    branch_req_4398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(186), ack => if_stmt_1576_branch_req_0); -- 
    -- CP-element group 187:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	882 
    -- CP-element group 187: 	883 
    -- CP-element group 187: 	885 
    -- CP-element group 187: 	886 
    -- CP-element group 187: 	888 
    -- CP-element group 187: 	889 
    -- CP-element group 187:  members (40) 
      -- CP-element group 187: 	 branch_block_stmt_655/merge_stmt_1582__exit__
      -- CP-element group 187: 	 branch_block_stmt_655/assign_stmt_1588__entry__
      -- CP-element group 187: 	 branch_block_stmt_655/assign_stmt_1588__exit__
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389
      -- CP-element group 187: 	 branch_block_stmt_655/if_stmt_1576_if_link/$exit
      -- CP-element group 187: 	 branch_block_stmt_655/if_stmt_1576_if_link/if_choice_transition
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xend338_ifx_xthen348
      -- CP-element group 187: 	 branch_block_stmt_655/assign_stmt_1588/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/assign_stmt_1588/$exit
      -- CP-element group 187: 	 branch_block_stmt_655/merge_stmt_1582_PhiReqMerge
      -- CP-element group 187: 	 branch_block_stmt_655/merge_stmt_1582_PhiAck/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/Update/cr
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xend338_ifx_xthen348_PhiReq/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xend338_ifx_xthen348_PhiReq/$exit
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/Update/cr
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/merge_stmt_1582_PhiAck/dummy
      -- CP-element group 187: 	 branch_block_stmt_655/merge_stmt_1582_PhiAck/$exit
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/Update/cr
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/$entry
      -- CP-element group 187: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/$entry
      -- 
    if_choice_transition_4403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1576_branch_ack_1, ack => zeropad3D_CP_2067_elements(187)); -- 
    rr_11370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(187), ack => type_cast_1680_inst_req_0); -- 
    cr_11375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(187), ack => type_cast_1680_inst_req_1); -- 
    cr_11398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(187), ack => type_cast_1672_inst_req_1); -- 
    rr_11393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(187), ack => type_cast_1672_inst_req_0); -- 
    cr_11352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(187), ack => type_cast_1684_inst_req_1); -- 
    rr_11347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(187), ack => type_cast_1684_inst_req_0); -- 
    -- CP-element group 188:  fork  transition  place  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	190 
    -- CP-element group 188: 	191 
    -- CP-element group 188: 	192 
    -- CP-element group 188: 	194 
    -- CP-element group 188: 	197 
    -- CP-element group 188: 	199 
    -- CP-element group 188: 	200 
    -- CP-element group 188: 	201 
    -- CP-element group 188: 	203 
    -- CP-element group 188:  members (54) 
      -- CP-element group 188: 	 branch_block_stmt_655/merge_stmt_1590__exit__
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661__entry__
      -- CP-element group 188: 	 branch_block_stmt_655/if_stmt_1576_else_link/$exit
      -- CP-element group 188: 	 branch_block_stmt_655/if_stmt_1576_else_link/else_choice_transition
      -- CP-element group 188: 	 branch_block_stmt_655/ifx_xend338_ifx_xelse353
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_update_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_update_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_word_address_calculated
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_root_address_calculated
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Sample/word_access_start/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Sample/word_access_start/word_0/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Sample/word_access_start/word_0/rr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/word_access_complete/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/word_access_complete/word_0/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/word_access_complete/word_0/cr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_update_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_update_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_update_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_update_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_word_address_calculated
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_root_address_calculated
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Sample/word_access_start/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Sample/word_access_start/word_0/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Sample/word_access_start/word_0/rr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/word_access_complete/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/word_access_complete/word_0/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/word_access_complete/word_0/cr
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_update_start_
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_Update/cr
      -- CP-element group 188: 	 branch_block_stmt_655/merge_stmt_1590_PhiReqMerge
      -- CP-element group 188: 	 branch_block_stmt_655/merge_stmt_1590_PhiAck/dummy
      -- CP-element group 188: 	 branch_block_stmt_655/merge_stmt_1590_PhiAck/$exit
      -- CP-element group 188: 	 branch_block_stmt_655/merge_stmt_1590_PhiAck/$entry
      -- CP-element group 188: 	 branch_block_stmt_655/ifx_xend338_ifx_xelse353_PhiReq/$exit
      -- CP-element group 188: 	 branch_block_stmt_655/ifx_xend338_ifx_xelse353_PhiReq/$entry
      -- 
    else_choice_transition_4407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1576_branch_ack_0, ack => zeropad3D_CP_2067_elements(188)); -- 
    rr_4423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => type_cast_1600_inst_req_0); -- 
    cr_4428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => type_cast_1600_inst_req_1); -- 
    rr_4445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => LOAD_col_high_1603_load_0_req_0); -- 
    cr_4456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => LOAD_col_high_1603_load_0_req_1); -- 
    cr_4475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => type_cast_1607_inst_req_1); -- 
    cr_4489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => type_cast_1621_inst_req_1); -- 
    cr_4503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => type_cast_1637_inst_req_1); -- 
    rr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => LOAD_row_high_1640_load_0_req_0); -- 
    cr_4531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => LOAD_row_high_1640_load_0_req_1); -- 
    cr_4550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(188), ack => type_cast_1644_inst_req_1); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_Sample/ra
      -- 
    ra_4424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1600_inst_ack_0, ack => zeropad3D_CP_2067_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	195 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1600_Update/ca
      -- 
    ca_4429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1600_inst_ack_1, ack => zeropad3D_CP_2067_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (5) 
      -- CP-element group 191: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Sample/word_access_start/$exit
      -- CP-element group 191: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Sample/word_access_start/word_0/$exit
      -- CP-element group 191: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Sample/word_access_start/word_0/ra
      -- 
    ra_4446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1603_load_0_ack_0, ack => zeropad3D_CP_2067_elements(191)); -- 
    -- CP-element group 192:  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	188 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (12) 
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/word_access_complete/$exit
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/word_access_complete/word_0/$exit
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/word_access_complete/word_0/ca
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/LOAD_col_high_1603_Merge/$entry
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/LOAD_col_high_1603_Merge/$exit
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/LOAD_col_high_1603_Merge/merge_req
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_col_high_1603_Update/LOAD_col_high_1603_Merge/merge_ack
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_Sample/rr
      -- 
    ca_4457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1603_load_0_ack_1, ack => zeropad3D_CP_2067_elements(192)); -- 
    rr_4470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(192), ack => type_cast_1607_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_Sample/ra
      -- 
    ra_4471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_0, ack => zeropad3D_CP_2067_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	188 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1607_Update/ca
      -- 
    ca_4476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_1, ack => zeropad3D_CP_2067_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	190 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_Sample/rr
      -- 
    rr_4484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(195), ack => type_cast_1621_inst_req_0); -- 
    zeropad3D_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(190) & zeropad3D_CP_2067_elements(194);
      gj_zeropad3D_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_Sample/ra
      -- 
    ra_4485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1621_inst_ack_0, ack => zeropad3D_CP_2067_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	188 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1621_Update/ca
      -- CP-element group 197: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_Sample/rr
      -- 
    ca_4490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1621_inst_ack_1, ack => zeropad3D_CP_2067_elements(197)); -- 
    rr_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(197), ack => type_cast_1637_inst_req_0); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_Sample/ra
      -- 
    ra_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1637_inst_ack_0, ack => zeropad3D_CP_2067_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	188 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	204 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1637_Update/ca
      -- 
    ca_4504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1637_inst_ack_1, ack => zeropad3D_CP_2067_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	188 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (5) 
      -- CP-element group 200: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Sample/word_access_start/$exit
      -- CP-element group 200: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Sample/word_access_start/word_0/$exit
      -- CP-element group 200: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Sample/word_access_start/word_0/ra
      -- 
    ra_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1640_load_0_ack_0, ack => zeropad3D_CP_2067_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	188 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (12) 
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/word_access_complete/$exit
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/word_access_complete/word_0/$exit
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/word_access_complete/word_0/ca
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/LOAD_row_high_1640_Merge/$entry
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/LOAD_row_high_1640_Merge/$exit
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/LOAD_row_high_1640_Merge/merge_req
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/LOAD_row_high_1640_Update/LOAD_row_high_1640_Merge/merge_ack
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_Sample/rr
      -- 
    ca_4532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1640_load_0_ack_1, ack => zeropad3D_CP_2067_elements(201)); -- 
    rr_4545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(201), ack => type_cast_1644_inst_req_0); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_Sample/ra
      -- 
    ra_4546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_0, ack => zeropad3D_CP_2067_elements(202)); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	188 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/type_cast_1644_Update/ca
      -- 
    ca_4551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_1, ack => zeropad3D_CP_2067_elements(203)); -- 
    -- CP-element group 204:  branch  join  transition  place  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	199 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (10) 
      -- CP-element group 204: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661__exit__
      -- CP-element group 204: 	 branch_block_stmt_655/if_stmt_1662__entry__
      -- CP-element group 204: 	 branch_block_stmt_655/assign_stmt_1596_to_assign_stmt_1661/$exit
      -- CP-element group 204: 	 branch_block_stmt_655/if_stmt_1662_dead_link/$entry
      -- CP-element group 204: 	 branch_block_stmt_655/if_stmt_1662_eval_test/$entry
      -- CP-element group 204: 	 branch_block_stmt_655/if_stmt_1662_eval_test/$exit
      -- CP-element group 204: 	 branch_block_stmt_655/if_stmt_1662_eval_test/branch_req
      -- CP-element group 204: 	 branch_block_stmt_655/R_cmp380_1663_place
      -- CP-element group 204: 	 branch_block_stmt_655/if_stmt_1662_if_link/$entry
      -- CP-element group 204: 	 branch_block_stmt_655/if_stmt_1662_else_link/$entry
      -- 
    branch_req_4559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(204), ack => if_stmt_1662_branch_req_0); -- 
    zeropad3D_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(199) & zeropad3D_CP_2067_elements(203);
      gj_zeropad3D_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  place  input  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	897 
    -- CP-element group 205: 	898 
    -- CP-element group 205: 	900 
    -- CP-element group 205: 	901 
    -- CP-element group 205:  members (20) 
      -- CP-element group 205: 	 branch_block_stmt_655/if_stmt_1662_if_link/$exit
      -- CP-element group 205: 	 branch_block_stmt_655/if_stmt_1662_if_link/if_choice_transition
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/Update/cr
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/Sample/rr
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/Update/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/Update/cr
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/Update/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/Sample/rr
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/$entry
      -- CP-element group 205: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/$entry
      -- 
    if_choice_transition_4564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1662_branch_ack_1, ack => zeropad3D_CP_2067_elements(205)); -- 
    cr_11454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(205), ack => type_cast_1694_inst_req_1); -- 
    rr_11449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(205), ack => type_cast_1694_inst_req_0); -- 
    cr_11431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(205), ack => type_cast_1698_inst_req_1); -- 
    rr_11426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(205), ack => type_cast_1698_inst_req_0); -- 
    -- CP-element group 206:  fork  transition  place  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	874 
    -- CP-element group 206: 	875 
    -- CP-element group 206: 	876 
    -- CP-element group 206: 	878 
    -- CP-element group 206: 	879 
    -- CP-element group 206:  members (22) 
      -- CP-element group 206: 	 branch_block_stmt_655/if_stmt_1662_else_link/$exit
      -- CP-element group 206: 	 branch_block_stmt_655/if_stmt_1662_else_link/else_choice_transition
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1681/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/Update/cr
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/Update/cr
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/Sample/rr
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/Sample/rr
      -- 
    else_choice_transition_4568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1662_branch_ack_0, ack => zeropad3D_CP_2067_elements(206)); -- 
    cr_11326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(206), ack => type_cast_1674_inst_req_1); -- 
    cr_11303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(206), ack => type_cast_1678_inst_req_1); -- 
    rr_11298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(206), ack => type_cast_1678_inst_req_0); -- 
    rr_11321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(206), ack => type_cast_1674_inst_req_0); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	906 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_Sample/ra
      -- 
    ra_4582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1702_inst_ack_0, ack => zeropad3D_CP_2067_elements(207)); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	906 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	227 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_Update/ca
      -- 
    ca_4587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1702_inst_ack_1, ack => zeropad3D_CP_2067_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	906 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Sample/word_access_start/$exit
      -- CP-element group 209: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Sample/word_access_start/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Sample/word_access_start/word_0/ra
      -- 
    ra_4604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1711_load_0_ack_0, ack => zeropad3D_CP_2067_elements(209)); -- 
    -- CP-element group 210:  transition  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	906 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	223 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/word_access_complete/$exit
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/word_access_complete/word_0/$exit
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/word_access_complete/word_0/ca
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/LOAD_pad_1711_Merge/$entry
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/LOAD_pad_1711_Merge/$exit
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/LOAD_pad_1711_Merge/merge_req
      -- CP-element group 210: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/LOAD_pad_1711_Merge/merge_ack
      -- 
    ca_4615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1711_load_0_ack_1, ack => zeropad3D_CP_2067_elements(210)); -- 
    rr_4769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(210), ack => type_cast_1741_inst_req_0); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	906 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (5) 
      -- CP-element group 211: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Sample/word_access_start/$exit
      -- CP-element group 211: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Sample/word_access_start/word_0/$exit
      -- CP-element group 211: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Sample/word_access_start/word_0/ra
      -- 
    ra_4637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1714_load_0_ack_0, ack => zeropad3D_CP_2067_elements(211)); -- 
    -- CP-element group 212:  transition  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	906 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (12) 
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/LOAD_depth_high_1714_Merge/merge_ack
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/LOAD_depth_high_1714_Merge/merge_req
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/LOAD_depth_high_1714_Merge/$exit
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/LOAD_depth_high_1714_Merge/$entry
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/word_access_complete/$exit
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/word_access_complete/word_0/$exit
      -- CP-element group 212: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/word_access_complete/word_0/ca
      -- 
    ca_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1714_load_0_ack_1, ack => zeropad3D_CP_2067_elements(212)); -- 
    rr_4727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(212), ack => type_cast_1724_inst_req_0); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	906 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Sample/word_access_start/word_0/ra
      -- CP-element group 213: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Sample/word_access_start/$exit
      -- CP-element group 213: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Sample/word_access_start/word_0/$exit
      -- CP-element group 213: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_sample_completed_
      -- 
    ra_4670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_1717_load_0_ack_0, ack => zeropad3D_CP_2067_elements(213)); -- 
    -- CP-element group 214:  fork  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	906 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	219 
    -- CP-element group 214: 	225 
    -- CP-element group 214:  members (15) 
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/LOAD_out_depth_high_1717_Merge/merge_ack
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/LOAD_out_depth_high_1717_Merge/merge_req
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/LOAD_out_depth_high_1717_Merge/$exit
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/LOAD_out_depth_high_1717_Merge/$entry
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/word_access_complete/word_0/ca
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/word_access_complete/word_0/$exit
      -- CP-element group 214: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/word_access_complete/$exit
      -- 
    ca_4681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_1717_load_0_ack_1, ack => zeropad3D_CP_2067_elements(214)); -- 
    rr_4741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(214), ack => type_cast_1728_inst_req_0); -- 
    rr_4783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(214), ack => type_cast_1745_inst_req_0); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	906 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (5) 
      -- CP-element group 215: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Sample/word_access_start/word_0/$exit
      -- CP-element group 215: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Sample/word_access_start/word_0/ra
      -- CP-element group 215: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Sample/word_access_start/$exit
      -- CP-element group 215: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_sample_completed_
      -- 
    ra_4703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_1720_load_0_ack_0, ack => zeropad3D_CP_2067_elements(215)); -- 
    -- CP-element group 216:  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	906 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	221 
    -- CP-element group 216:  members (12) 
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/LOAD_out_col_high_1720_Merge/$exit
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/LOAD_out_col_high_1720_Merge/merge_req
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/LOAD_out_col_high_1720_Merge/merge_ack
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/word_access_complete/$exit
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/word_access_complete/word_0/$exit
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_Sample/rr
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/LOAD_out_col_high_1720_Merge/$entry
      -- CP-element group 216: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/word_access_complete/word_0/ca
      -- 
    ca_4714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_1720_load_0_ack_1, ack => zeropad3D_CP_2067_elements(216)); -- 
    rr_4755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(216), ack => type_cast_1732_inst_req_0); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_sample_completed_
      -- 
    ra_4728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1724_inst_ack_0, ack => zeropad3D_CP_2067_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	906 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	227 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_update_completed_
      -- 
    ca_4733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1724_inst_ack_1, ack => zeropad3D_CP_2067_elements(218)); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	214 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_Sample/ra
      -- CP-element group 219: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_sample_completed_
      -- 
    ra_4742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1728_inst_ack_0, ack => zeropad3D_CP_2067_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	906 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	227 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_Update/ca
      -- CP-element group 220: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_update_completed_
      -- 
    ca_4747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1728_inst_ack_1, ack => zeropad3D_CP_2067_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	216 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_Sample/ra
      -- CP-element group 221: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_sample_completed_
      -- 
    ra_4756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1732_inst_ack_0, ack => zeropad3D_CP_2067_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	906 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	227 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_Update/ca
      -- CP-element group 222: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_update_completed_
      -- 
    ca_4761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1732_inst_ack_1, ack => zeropad3D_CP_2067_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	210 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_Sample/ra
      -- 
    ra_4770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1741_inst_ack_0, ack => zeropad3D_CP_2067_elements(223)); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	906 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	227 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_Update/ca
      -- 
    ca_4775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1741_inst_ack_1, ack => zeropad3D_CP_2067_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	214 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_Sample/ra
      -- CP-element group 225: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_Sample/$exit
      -- 
    ra_4784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1745_inst_ack_0, ack => zeropad3D_CP_2067_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	906 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_Update/ca
      -- CP-element group 226: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_update_completed_
      -- 
    ca_4789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1745_inst_ack_1, ack => zeropad3D_CP_2067_elements(226)); -- 
    -- CP-element group 227:  join  fork  transition  place  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	208 
    -- CP-element group 227: 	218 
    -- CP-element group 227: 	220 
    -- CP-element group 227: 	222 
    -- CP-element group 227: 	224 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	917 
    -- CP-element group 227: 	918 
    -- CP-element group 227: 	919 
    -- CP-element group 227: 	921 
    -- CP-element group 227:  members (16) 
      -- CP-element group 227: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787__exit__
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450
      -- CP-element group 227: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/$exit
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Update/cr
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Sample/rr
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1803/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1790/$entry
      -- CP-element group 227: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/$entry
      -- 
    cr_11566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(227), ack => type_cast_1800_inst_req_1); -- 
    rr_11561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(227), ack => type_cast_1800_inst_req_0); -- 
    zeropad3D_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(208) & zeropad3D_CP_2067_elements(218) & zeropad3D_CP_2067_elements(220) & zeropad3D_CP_2067_elements(222) & zeropad3D_CP_2067_elements(224) & zeropad3D_CP_2067_elements(226);
      gj_zeropad3D_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	927 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_Sample/ra
      -- CP-element group 228: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_sample_completed_
      -- 
    ra_4801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1814_inst_ack_0, ack => zeropad3D_CP_2067_elements(228)); -- 
    -- CP-element group 229:  branch  transition  place  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	927 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822__exit__
      -- CP-element group 229: 	 branch_block_stmt_655/if_stmt_1823__entry__
      -- CP-element group 229: 	 branch_block_stmt_655/if_stmt_1823_dead_link/$entry
      -- CP-element group 229: 	 branch_block_stmt_655/if_stmt_1823_eval_test/$entry
      -- CP-element group 229: 	 branch_block_stmt_655/if_stmt_1823_eval_test/$exit
      -- CP-element group 229: 	 branch_block_stmt_655/if_stmt_1823_eval_test/branch_req
      -- CP-element group 229: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_Update/ca
      -- CP-element group 229: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/$exit
      -- CP-element group 229: 	 branch_block_stmt_655/if_stmt_1823_else_link/$entry
      -- CP-element group 229: 	 branch_block_stmt_655/R_cmp455_1824_place
      -- CP-element group 229: 	 branch_block_stmt_655/if_stmt_1823_if_link/$entry
      -- 
    ca_4806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1814_inst_ack_1, ack => zeropad3D_CP_2067_elements(229)); -- 
    branch_req_4814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(229), ack => if_stmt_1823_branch_req_0); -- 
    -- CP-element group 230:  transition  place  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	928 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_655/whilex_xbody450_ifx_xthen486
      -- CP-element group 230: 	 branch_block_stmt_655/if_stmt_1823_if_link/if_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_655/if_stmt_1823_if_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_655/whilex_xbody450_ifx_xthen486_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_655/whilex_xbody450_ifx_xthen486_PhiReq/$exit
      -- 
    if_choice_transition_4819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1823_branch_ack_1, ack => zeropad3D_CP_2067_elements(230)); -- 
    -- CP-element group 231:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231: 	233 
    -- CP-element group 231: 	235 
    -- CP-element group 231:  members (27) 
      -- CP-element group 231: 	 branch_block_stmt_655/merge_stmt_1829__exit__
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854__entry__
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_root_address_calculated
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/word_access_complete/word_0/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/word_access_complete/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Sample/word_access_start/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/word_access_complete/word_0/cr
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Sample/word_access_start/word_0/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Sample/word_access_start/word_0/rr
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_word_address_calculated
      -- CP-element group 231: 	 branch_block_stmt_655/whilex_xbody450_lorx_xlhsx_xfalse457
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_update_start_
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_update_start_
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/if_stmt_1823_else_link/else_choice_transition
      -- CP-element group 231: 	 branch_block_stmt_655/if_stmt_1823_else_link/$exit
      -- CP-element group 231: 	 branch_block_stmt_655/merge_stmt_1829_PhiReqMerge
      -- CP-element group 231: 	 branch_block_stmt_655/whilex_xbody450_lorx_xlhsx_xfalse457_PhiReq/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/whilex_xbody450_lorx_xlhsx_xfalse457_PhiReq/$exit
      -- CP-element group 231: 	 branch_block_stmt_655/merge_stmt_1829_PhiAck/$entry
      -- CP-element group 231: 	 branch_block_stmt_655/merge_stmt_1829_PhiAck/$exit
      -- CP-element group 231: 	 branch_block_stmt_655/merge_stmt_1829_PhiAck/dummy
      -- 
    else_choice_transition_4823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1823_branch_ack_0, ack => zeropad3D_CP_2067_elements(231)); -- 
    cr_4874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(231), ack => type_cast_1835_inst_req_1); -- 
    cr_4855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(231), ack => LOAD_row_high_1831_load_0_req_1); -- 
    rr_4844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(231), ack => LOAD_row_high_1831_load_0_req_0); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (5) 
      -- CP-element group 232: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Sample/word_access_start/$exit
      -- CP-element group 232: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Sample/word_access_start/word_0/$exit
      -- CP-element group 232: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Sample/word_access_start/word_0/ra
      -- CP-element group 232: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_sample_completed_
      -- 
    ra_4845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1831_load_0_ack_0, ack => zeropad3D_CP_2067_elements(232)); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (12) 
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/word_access_complete/word_0/ca
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/word_access_complete/word_0/$exit
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/word_access_complete/$exit
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_Sample/rr
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/LOAD_row_high_1831_Merge/merge_ack
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/LOAD_row_high_1831_Merge/merge_req
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/LOAD_row_high_1831_Merge/$exit
      -- CP-element group 233: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/LOAD_row_high_1831_Update/LOAD_row_high_1831_Merge/$entry
      -- 
    ca_4856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1831_load_0_ack_1, ack => zeropad3D_CP_2067_elements(233)); -- 
    rr_4869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(233), ack => type_cast_1835_inst_req_0); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_Sample/ra
      -- CP-element group 234: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_sample_completed_
      -- 
    ra_4870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_0, ack => zeropad3D_CP_2067_elements(234)); -- 
    -- CP-element group 235:  branch  transition  place  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	231 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (13) 
      -- CP-element group 235: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854__exit__
      -- CP-element group 235: 	 branch_block_stmt_655/if_stmt_1855__entry__
      -- CP-element group 235: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_Update/ca
      -- CP-element group 235: 	 branch_block_stmt_655/if_stmt_1855_dead_link/$entry
      -- CP-element group 235: 	 branch_block_stmt_655/if_stmt_1855_eval_test/$entry
      -- CP-element group 235: 	 branch_block_stmt_655/if_stmt_1855_eval_test/$exit
      -- CP-element group 235: 	 branch_block_stmt_655/R_cmp466_1856_place
      -- CP-element group 235: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/type_cast_1835_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_655/assign_stmt_1832_to_assign_stmt_1854/$exit
      -- CP-element group 235: 	 branch_block_stmt_655/if_stmt_1855_else_link/$entry
      -- CP-element group 235: 	 branch_block_stmt_655/if_stmt_1855_if_link/$entry
      -- CP-element group 235: 	 branch_block_stmt_655/if_stmt_1855_eval_test/branch_req
      -- 
    ca_4875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_1, ack => zeropad3D_CP_2067_elements(235)); -- 
    branch_req_4883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(235), ack => if_stmt_1855_branch_req_0); -- 
    -- CP-element group 236:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236: 	239 
    -- CP-element group 236:  members (18) 
      -- CP-element group 236: 	 branch_block_stmt_655/merge_stmt_1861__exit__
      -- CP-element group 236: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873__entry__
      -- CP-element group 236: 	 branch_block_stmt_655/lorx_xlhsx_xfalse457_lorx_xlhsx_xfalse468
      -- CP-element group 236: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/$entry
      -- CP-element group 236: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_655/if_stmt_1855_if_link/if_choice_transition
      -- CP-element group 236: 	 branch_block_stmt_655/if_stmt_1855_if_link/$exit
      -- CP-element group 236: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_update_start_
      -- CP-element group 236: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_Sample/rr
      -- CP-element group 236: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_Update/$entry
      -- CP-element group 236: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_Update/cr
      -- CP-element group 236: 	 branch_block_stmt_655/merge_stmt_1861_PhiReqMerge
      -- CP-element group 236: 	 branch_block_stmt_655/lorx_xlhsx_xfalse457_lorx_xlhsx_xfalse468_PhiReq/$entry
      -- CP-element group 236: 	 branch_block_stmt_655/lorx_xlhsx_xfalse457_lorx_xlhsx_xfalse468_PhiReq/$exit
      -- CP-element group 236: 	 branch_block_stmt_655/merge_stmt_1861_PhiAck/$entry
      -- CP-element group 236: 	 branch_block_stmt_655/merge_stmt_1861_PhiAck/$exit
      -- CP-element group 236: 	 branch_block_stmt_655/merge_stmt_1861_PhiAck/dummy
      -- 
    if_choice_transition_4888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1855_branch_ack_1, ack => zeropad3D_CP_2067_elements(236)); -- 
    rr_4905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(236), ack => type_cast_1865_inst_req_0); -- 
    cr_4910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(236), ack => type_cast_1865_inst_req_1); -- 
    -- CP-element group 237:  transition  place  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	928 
    -- CP-element group 237:  members (5) 
      -- CP-element group 237: 	 branch_block_stmt_655/lorx_xlhsx_xfalse457_ifx_xthen486
      -- CP-element group 237: 	 branch_block_stmt_655/if_stmt_1855_else_link/else_choice_transition
      -- CP-element group 237: 	 branch_block_stmt_655/if_stmt_1855_else_link/$exit
      -- CP-element group 237: 	 branch_block_stmt_655/lorx_xlhsx_xfalse457_ifx_xthen486_PhiReq/$entry
      -- CP-element group 237: 	 branch_block_stmt_655/lorx_xlhsx_xfalse457_ifx_xthen486_PhiReq/$exit
      -- 
    else_choice_transition_4892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1855_branch_ack_0, ack => zeropad3D_CP_2067_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_sample_completed_
      -- CP-element group 238: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_Sample/ra
      -- 
    ra_4906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_0, ack => zeropad3D_CP_2067_elements(238)); -- 
    -- CP-element group 239:  branch  transition  place  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	236 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (13) 
      -- CP-element group 239: 	 branch_block_stmt_655/if_stmt_1874__entry__
      -- CP-element group 239: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873__exit__
      -- CP-element group 239: 	 branch_block_stmt_655/R_cmp473_1875_place
      -- CP-element group 239: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/$exit
      -- CP-element group 239: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_655/assign_stmt_1866_to_assign_stmt_1873/type_cast_1865_Update/ca
      -- CP-element group 239: 	 branch_block_stmt_655/if_stmt_1874_dead_link/$entry
      -- CP-element group 239: 	 branch_block_stmt_655/if_stmt_1874_eval_test/$entry
      -- CP-element group 239: 	 branch_block_stmt_655/if_stmt_1874_eval_test/$exit
      -- CP-element group 239: 	 branch_block_stmt_655/if_stmt_1874_eval_test/branch_req
      -- CP-element group 239: 	 branch_block_stmt_655/if_stmt_1874_if_link/$entry
      -- CP-element group 239: 	 branch_block_stmt_655/if_stmt_1874_else_link/$entry
      -- 
    ca_4911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_1, ack => zeropad3D_CP_2067_elements(239)); -- 
    branch_req_4919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(239), ack => if_stmt_1874_branch_req_0); -- 
    -- CP-element group 240:  transition  place  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	928 
    -- CP-element group 240:  members (5) 
      -- CP-element group 240: 	 branch_block_stmt_655/lorx_xlhsx_xfalse468_ifx_xthen486
      -- CP-element group 240: 	 branch_block_stmt_655/if_stmt_1874_if_link/$exit
      -- CP-element group 240: 	 branch_block_stmt_655/if_stmt_1874_if_link/if_choice_transition
      -- CP-element group 240: 	 branch_block_stmt_655/lorx_xlhsx_xfalse468_ifx_xthen486_PhiReq/$entry
      -- CP-element group 240: 	 branch_block_stmt_655/lorx_xlhsx_xfalse468_ifx_xthen486_PhiReq/$exit
      -- 
    if_choice_transition_4924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1874_branch_ack_1, ack => zeropad3D_CP_2067_elements(240)); -- 
    -- CP-element group 241:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241: 	243 
    -- CP-element group 241: 	245 
    -- CP-element group 241:  members (27) 
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905__entry__
      -- CP-element group 241: 	 branch_block_stmt_655/merge_stmt_1880__exit__
      -- CP-element group 241: 	 branch_block_stmt_655/lorx_xlhsx_xfalse468_lorx_xlhsx_xfalse475
      -- CP-element group 241: 	 branch_block_stmt_655/if_stmt_1874_else_link/$exit
      -- CP-element group 241: 	 branch_block_stmt_655/if_stmt_1874_else_link/else_choice_transition
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_update_start_
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_word_address_calculated
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_root_address_calculated
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Sample/word_access_start/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Sample/word_access_start/word_0/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Sample/word_access_start/word_0/rr
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/word_access_complete/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/word_access_complete/word_0/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/word_access_complete/word_0/cr
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_update_start_
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_Update/cr
      -- CP-element group 241: 	 branch_block_stmt_655/merge_stmt_1880_PhiReqMerge
      -- CP-element group 241: 	 branch_block_stmt_655/lorx_xlhsx_xfalse468_lorx_xlhsx_xfalse475_PhiReq/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/lorx_xlhsx_xfalse468_lorx_xlhsx_xfalse475_PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_655/merge_stmt_1880_PhiAck/$entry
      -- CP-element group 241: 	 branch_block_stmt_655/merge_stmt_1880_PhiAck/$exit
      -- CP-element group 241: 	 branch_block_stmt_655/merge_stmt_1880_PhiAck/dummy
      -- 
    else_choice_transition_4928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1874_branch_ack_0, ack => zeropad3D_CP_2067_elements(241)); -- 
    rr_4949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(241), ack => LOAD_col_high_1882_load_0_req_0); -- 
    cr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(241), ack => LOAD_col_high_1882_load_0_req_1); -- 
    cr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(241), ack => type_cast_1886_inst_req_1); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (5) 
      -- CP-element group 242: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_sample_completed_
      -- CP-element group 242: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Sample/word_access_start/$exit
      -- CP-element group 242: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Sample/word_access_start/word_0/$exit
      -- CP-element group 242: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Sample/word_access_start/word_0/ra
      -- 
    ra_4950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1882_load_0_ack_0, ack => zeropad3D_CP_2067_elements(242)); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (12) 
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/word_access_complete/$exit
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/word_access_complete/word_0/$exit
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/word_access_complete/word_0/ca
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/LOAD_col_high_1882_Merge/$entry
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/LOAD_col_high_1882_Merge/$exit
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/LOAD_col_high_1882_Merge/merge_req
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/LOAD_col_high_1882_Update/LOAD_col_high_1882_Merge/merge_ack
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_Sample/rr
      -- 
    ca_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1882_load_0_ack_1, ack => zeropad3D_CP_2067_elements(243)); -- 
    rr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(243), ack => type_cast_1886_inst_req_0); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_Sample/ra
      -- 
    ra_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1886_inst_ack_0, ack => zeropad3D_CP_2067_elements(244)); -- 
    -- CP-element group 245:  branch  transition  place  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	241 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (13) 
      -- CP-element group 245: 	 branch_block_stmt_655/if_stmt_1906__entry__
      -- CP-element group 245: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905__exit__
      -- CP-element group 245: 	 branch_block_stmt_655/R_cmp484_1907_place
      -- CP-element group 245: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/$exit
      -- CP-element group 245: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_655/assign_stmt_1883_to_assign_stmt_1905/type_cast_1886_Update/ca
      -- CP-element group 245: 	 branch_block_stmt_655/if_stmt_1906_dead_link/$entry
      -- CP-element group 245: 	 branch_block_stmt_655/if_stmt_1906_eval_test/$entry
      -- CP-element group 245: 	 branch_block_stmt_655/if_stmt_1906_eval_test/$exit
      -- CP-element group 245: 	 branch_block_stmt_655/if_stmt_1906_eval_test/branch_req
      -- CP-element group 245: 	 branch_block_stmt_655/if_stmt_1906_if_link/$entry
      -- CP-element group 245: 	 branch_block_stmt_655/if_stmt_1906_else_link/$entry
      -- 
    ca_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1886_inst_ack_1, ack => zeropad3D_CP_2067_elements(245)); -- 
    branch_req_4988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(245), ack => if_stmt_1906_branch_req_0); -- 
    -- CP-element group 246:  fork  transition  place  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	262 
    -- CP-element group 246: 	263 
    -- CP-element group 246: 	265 
    -- CP-element group 246: 	267 
    -- CP-element group 246: 	269 
    -- CP-element group 246: 	271 
    -- CP-element group 246: 	273 
    -- CP-element group 246: 	275 
    -- CP-element group 246: 	277 
    -- CP-element group 246: 	280 
    -- CP-element group 246:  members (46) 
      -- CP-element group 246: 	 branch_block_stmt_655/merge_stmt_1970__exit__
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075__entry__
      -- CP-element group 246: 	 branch_block_stmt_655/lorx_xlhsx_xfalse475_ifx_xelse507
      -- CP-element group 246: 	 branch_block_stmt_655/if_stmt_1906_if_link/$exit
      -- CP-element group 246: 	 branch_block_stmt_655/if_stmt_1906_if_link/if_choice_transition
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_update_start_
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_Sample/rr
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_Update/cr
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_update_start_
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_Update/cr
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_update_start_
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_update_start
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_Update/req
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_complete/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_complete/req
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_update_start_
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/word_access_complete/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/word_access_complete/word_0/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/word_access_complete/word_0/cr
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_update_start_
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_Update/cr
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_update_start_
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_update_start
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_Update/req
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_complete/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_complete/req
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_update_start_
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Update/word_access_complete/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Update/word_access_complete/word_0/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Update/word_access_complete/word_0/cr
      -- CP-element group 246: 	 branch_block_stmt_655/merge_stmt_1970_PhiReqMerge
      -- CP-element group 246: 	 branch_block_stmt_655/lorx_xlhsx_xfalse475_ifx_xelse507_PhiReq/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/lorx_xlhsx_xfalse475_ifx_xelse507_PhiReq/$exit
      -- CP-element group 246: 	 branch_block_stmt_655/merge_stmt_1970_PhiAck/$entry
      -- CP-element group 246: 	 branch_block_stmt_655/merge_stmt_1970_PhiAck/$exit
      -- CP-element group 246: 	 branch_block_stmt_655/merge_stmt_1970_PhiAck/dummy
      -- 
    if_choice_transition_4993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1906_branch_ack_1, ack => zeropad3D_CP_2067_elements(246)); -- 
    rr_5151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => type_cast_1974_inst_req_0); -- 
    cr_5156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => type_cast_1974_inst_req_1); -- 
    cr_5170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => type_cast_2038_inst_req_1); -- 
    req_5201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => array_obj_ref_2044_index_offset_req_1); -- 
    req_5216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => addr_of_2045_final_reg_req_1); -- 
    cr_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => ptr_deref_2049_load_0_req_1); -- 
    cr_5280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => type_cast_2063_inst_req_1); -- 
    req_5311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => array_obj_ref_2069_index_offset_req_1); -- 
    req_5326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => addr_of_2070_final_reg_req_1); -- 
    cr_5376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(246), ack => ptr_deref_2073_store_0_req_1); -- 
    -- CP-element group 247:  transition  place  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	928 
    -- CP-element group 247:  members (5) 
      -- CP-element group 247: 	 branch_block_stmt_655/lorx_xlhsx_xfalse475_ifx_xthen486
      -- CP-element group 247: 	 branch_block_stmt_655/if_stmt_1906_else_link/$exit
      -- CP-element group 247: 	 branch_block_stmt_655/if_stmt_1906_else_link/else_choice_transition
      -- CP-element group 247: 	 branch_block_stmt_655/lorx_xlhsx_xfalse475_ifx_xthen486_PhiReq/$entry
      -- CP-element group 247: 	 branch_block_stmt_655/lorx_xlhsx_xfalse475_ifx_xthen486_PhiReq/$exit
      -- 
    else_choice_transition_4997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1906_branch_ack_0, ack => zeropad3D_CP_2067_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	928 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_Sample/ra
      -- 
    ra_5011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1916_inst_ack_0, ack => zeropad3D_CP_2067_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	928 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	252 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_Update/ca
      -- 
    ca_5016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1916_inst_ack_1, ack => zeropad3D_CP_2067_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	928 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_Sample/ra
      -- 
    ra_5025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1921_inst_ack_0, ack => zeropad3D_CP_2067_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	928 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_Update/ca
      -- 
    ca_5030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1921_inst_ack_1, ack => zeropad3D_CP_2067_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	249 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_Sample/rr
      -- 
    rr_5038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(252), ack => type_cast_1955_inst_req_0); -- 
    zeropad3D_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(249) & zeropad3D_CP_2067_elements(251);
      gj_zeropad3D_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_Sample/ra
      -- 
    ra_5039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1955_inst_ack_0, ack => zeropad3D_CP_2067_elements(253)); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	928 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (16) 
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_Update/ca
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_resized_1
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_scaled_1
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_computed_1
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_resize_1/$entry
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_resize_1/$exit
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_resize_1/index_resize_req
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_resize_1/index_resize_ack
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_scale_1/$entry
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_scale_1/$exit
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_scale_1/scale_rename_req
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_index_scale_1/scale_rename_ack
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_Sample/req
      -- 
    ca_5044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1955_inst_ack_1, ack => zeropad3D_CP_2067_elements(254)); -- 
    req_5069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(254), ack => array_obj_ref_1961_index_offset_req_0); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	261 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_sample_complete
      -- CP-element group 255: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_Sample/ack
      -- 
    ack_5070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1961_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(255)); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	928 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (11) 
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_root_address_calculated
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_offset_calculated
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_base_plus_offset/$entry
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_base_plus_offset/$exit
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_base_plus_offset/sum_rename_req
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_base_plus_offset/sum_rename_ack
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_request/$entry
      -- CP-element group 256: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_request/req
      -- 
    ack_5075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1961_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(256)); -- 
    req_5084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(256), ack => addr_of_1962_final_reg_req_0); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_request/$exit
      -- CP-element group 257: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_request/ack
      -- 
    ack_5085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1962_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(257)); -- 
    -- CP-element group 258:  join  fork  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	928 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (28) 
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_complete/$exit
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_complete/ack
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_address_calculated
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_word_address_calculated
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_root_address_calculated
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_address_resized
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_addr_resize/$entry
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_addr_resize/$exit
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_addr_resize/base_resize_req
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_addr_resize/base_resize_ack
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_plus_offset/$entry
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_plus_offset/$exit
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_plus_offset/sum_rename_req
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_base_plus_offset/sum_rename_ack
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_word_addrgen/$entry
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_word_addrgen/$exit
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_word_addrgen/root_register_req
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_word_addrgen/root_register_ack
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/ptr_deref_1965_Split/$entry
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/ptr_deref_1965_Split/$exit
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/ptr_deref_1965_Split/split_req
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/ptr_deref_1965_Split/split_ack
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/word_access_start/$entry
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/word_access_start/word_0/$entry
      -- CP-element group 258: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/word_access_start/word_0/rr
      -- 
    ack_5090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1962_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(258)); -- 
    rr_5128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(258), ack => ptr_deref_1965_store_0_req_0); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259:  members (5) 
      -- CP-element group 259: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/word_access_start/$exit
      -- CP-element group 259: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/word_access_start/word_0/$exit
      -- CP-element group 259: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Sample/word_access_start/word_0/ra
      -- 
    ra_5129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1965_store_0_ack_0, ack => zeropad3D_CP_2067_elements(259)); -- 
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	928 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (5) 
      -- CP-element group 260: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Update/word_access_complete/$exit
      -- CP-element group 260: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Update/word_access_complete/word_0/$exit
      -- CP-element group 260: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Update/word_access_complete/word_0/ca
      -- 
    ca_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1965_store_0_ack_1, ack => zeropad3D_CP_2067_elements(260)); -- 
    -- CP-element group 261:  join  transition  place  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	255 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	929 
    -- CP-element group 261:  members (5) 
      -- CP-element group 261: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968__exit__
      -- CP-element group 261: 	 branch_block_stmt_655/ifx_xthen486_ifx_xend555
      -- CP-element group 261: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/$exit
      -- CP-element group 261: 	 branch_block_stmt_655/ifx_xthen486_ifx_xend555_PhiReq/$entry
      -- CP-element group 261: 	 branch_block_stmt_655/ifx_xthen486_ifx_xend555_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(255) & zeropad3D_CP_2067_elements(260);
      gj_zeropad3D_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	246 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_Sample/ra
      -- 
    ra_5152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1974_inst_ack_0, ack => zeropad3D_CP_2067_elements(262)); -- 
    -- CP-element group 263:  fork  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	246 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263: 	272 
    -- CP-element group 263:  members (9) 
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_1974_Update/ca
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_Sample/rr
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_Sample/rr
      -- 
    ca_5157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1974_inst_ack_1, ack => zeropad3D_CP_2067_elements(263)); -- 
    rr_5165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(263), ack => type_cast_2038_inst_req_0); -- 
    rr_5275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(263), ack => type_cast_2063_inst_req_0); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_Sample/ra
      -- 
    ra_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_0, ack => zeropad3D_CP_2067_elements(264)); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	246 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (16) 
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2038_Update/ca
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_resized_1
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_scaled_1
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_computed_1
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_resize_1/$entry
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_resize_1/$exit
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_resize_1/index_resize_req
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_resize_1/index_resize_ack
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_scale_1/$entry
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_scale_1/$exit
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_scale_1/scale_rename_req
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_index_scale_1/scale_rename_ack
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_Sample/req
      -- 
    ca_5171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_1, ack => zeropad3D_CP_2067_elements(265)); -- 
    req_5196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(265), ack => array_obj_ref_2044_index_offset_req_0); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	281 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_sample_complete
      -- CP-element group 266: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_Sample/ack
      -- 
    ack_5197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2044_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(266)); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	246 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (11) 
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_root_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_offset_calculated
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_final_index_sum_regn_Update/ack
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_base_plus_offset/$entry
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_base_plus_offset/$exit
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_base_plus_offset/sum_rename_req
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2044_base_plus_offset/sum_rename_ack
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_request/$entry
      -- CP-element group 267: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_request/req
      -- 
    ack_5202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2044_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(267)); -- 
    req_5211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(267), ack => addr_of_2045_final_reg_req_0); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_request/$exit
      -- CP-element group 268: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_request/ack
      -- 
    ack_5212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2045_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(268)); -- 
    -- CP-element group 269:  join  fork  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	246 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (24) 
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_complete/$exit
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2045_complete/ack
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_word_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_root_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_address_resized
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_addr_resize/$entry
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_addr_resize/$exit
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_addr_resize/base_resize_req
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_addr_resize/base_resize_ack
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_plus_offset/$entry
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_plus_offset/$exit
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_plus_offset/sum_rename_req
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_base_plus_offset/sum_rename_ack
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_word_addrgen/$entry
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_word_addrgen/$exit
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_word_addrgen/root_register_req
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_word_addrgen/root_register_ack
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Sample/word_access_start/$entry
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Sample/word_access_start/word_0/$entry
      -- CP-element group 269: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Sample/word_access_start/word_0/rr
      -- 
    ack_5217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2045_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(269)); -- 
    rr_5250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(269), ack => ptr_deref_2049_load_0_req_0); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (5) 
      -- CP-element group 270: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Sample/word_access_start/$exit
      -- CP-element group 270: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Sample/word_access_start/word_0/$exit
      -- CP-element group 270: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Sample/word_access_start/word_0/ra
      -- 
    ra_5251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2049_load_0_ack_0, ack => zeropad3D_CP_2067_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	246 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	278 
    -- CP-element group 271:  members (9) 
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/word_access_complete/$exit
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/word_access_complete/word_0/$exit
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/word_access_complete/word_0/ca
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/ptr_deref_2049_Merge/$entry
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/ptr_deref_2049_Merge/$exit
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/ptr_deref_2049_Merge/merge_req
      -- CP-element group 271: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2049_Update/ptr_deref_2049_Merge/merge_ack
      -- 
    ca_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2049_load_0_ack_1, ack => zeropad3D_CP_2067_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	263 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_Sample/ra
      -- 
    ra_5276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2063_inst_ack_0, ack => zeropad3D_CP_2067_elements(272)); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	246 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (16) 
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/type_cast_2063_Update/ca
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_resized_1
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_scaled_1
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_computed_1
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_resize_1/$entry
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_resize_1/$exit
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_resize_1/index_resize_req
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_resize_1/index_resize_ack
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_scale_1/$entry
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_scale_1/$exit
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_scale_1/scale_rename_req
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_index_scale_1/scale_rename_ack
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_Sample/req
      -- 
    ca_5281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2063_inst_ack_1, ack => zeropad3D_CP_2067_elements(273)); -- 
    req_5306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(273), ack => array_obj_ref_2069_index_offset_req_0); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	281 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_sample_complete
      -- CP-element group 274: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_Sample/ack
      -- 
    ack_5307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2069_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(274)); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	246 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (11) 
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_root_address_calculated
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_offset_calculated
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_final_index_sum_regn_Update/ack
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_base_plus_offset/$entry
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_base_plus_offset/$exit
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_base_plus_offset/sum_rename_req
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/array_obj_ref_2069_base_plus_offset/sum_rename_ack
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_request/$entry
      -- CP-element group 275: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_request/req
      -- 
    ack_5312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2069_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(275)); -- 
    req_5321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(275), ack => addr_of_2070_final_reg_req_0); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_request/$exit
      -- CP-element group 276: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_request/ack
      -- 
    ack_5322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2070_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(276)); -- 
    -- CP-element group 277:  fork  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	246 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (19) 
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_complete/$exit
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/addr_of_2070_complete/ack
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_address_calculated
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_word_address_calculated
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_root_address_calculated
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_address_resized
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_addr_resize/$entry
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_addr_resize/$exit
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_addr_resize/base_resize_req
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_addr_resize/base_resize_ack
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_plus_offset/$entry
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_plus_offset/$exit
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_plus_offset/sum_rename_req
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_base_plus_offset/sum_rename_ack
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_word_addrgen/$entry
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_word_addrgen/$exit
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_word_addrgen/root_register_req
      -- CP-element group 277: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_word_addrgen/root_register_ack
      -- 
    ack_5327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2070_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(277)); -- 
    -- CP-element group 278:  join  transition  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	271 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (9) 
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/ptr_deref_2073_Split/$entry
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/ptr_deref_2073_Split/$exit
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/ptr_deref_2073_Split/split_req
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/ptr_deref_2073_Split/split_ack
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/word_access_start/$entry
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/word_access_start/word_0/$entry
      -- CP-element group 278: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/word_access_start/word_0/rr
      -- 
    rr_5365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(278), ack => ptr_deref_2073_store_0_req_0); -- 
    zeropad3D_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(271) & zeropad3D_CP_2067_elements(277);
      gj_zeropad3D_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (5) 
      -- CP-element group 279: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/word_access_start/$exit
      -- CP-element group 279: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/word_access_start/word_0/$exit
      -- CP-element group 279: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Sample/word_access_start/word_0/ra
      -- 
    ra_5366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2073_store_0_ack_0, ack => zeropad3D_CP_2067_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	246 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (5) 
      -- CP-element group 280: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Update/word_access_complete/$exit
      -- CP-element group 280: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Update/word_access_complete/word_0/$exit
      -- CP-element group 280: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/ptr_deref_2073_Update/word_access_complete/word_0/ca
      -- 
    ca_5377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2073_store_0_ack_1, ack => zeropad3D_CP_2067_elements(280)); -- 
    -- CP-element group 281:  join  transition  place  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	266 
    -- CP-element group 281: 	274 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	929 
    -- CP-element group 281:  members (5) 
      -- CP-element group 281: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075__exit__
      -- CP-element group 281: 	 branch_block_stmt_655/ifx_xelse507_ifx_xend555
      -- CP-element group 281: 	 branch_block_stmt_655/assign_stmt_1975_to_assign_stmt_2075/$exit
      -- CP-element group 281: 	 branch_block_stmt_655/ifx_xelse507_ifx_xend555_PhiReq/$entry
      -- CP-element group 281: 	 branch_block_stmt_655/ifx_xelse507_ifx_xend555_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(266) & zeropad3D_CP_2067_elements(274) & zeropad3D_CP_2067_elements(280);
      gj_zeropad3D_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	929 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_sample_completed_
      -- CP-element group 282: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_Sample/ra
      -- 
    ra_5389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2081_inst_ack_0, ack => zeropad3D_CP_2067_elements(282)); -- 
    -- CP-element group 283:  branch  transition  place  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	929 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (13) 
      -- CP-element group 283: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095__exit__
      -- CP-element group 283: 	 branch_block_stmt_655/if_stmt_2096__entry__
      -- CP-element group 283: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/$exit
      -- CP-element group 283: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_update_completed_
      -- CP-element group 283: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_Update/ca
      -- CP-element group 283: 	 branch_block_stmt_655/if_stmt_2096_dead_link/$entry
      -- CP-element group 283: 	 branch_block_stmt_655/if_stmt_2096_eval_test/$entry
      -- CP-element group 283: 	 branch_block_stmt_655/if_stmt_2096_eval_test/$exit
      -- CP-element group 283: 	 branch_block_stmt_655/if_stmt_2096_eval_test/branch_req
      -- CP-element group 283: 	 branch_block_stmt_655/R_cmp563_2097_place
      -- CP-element group 283: 	 branch_block_stmt_655/if_stmt_2096_if_link/$entry
      -- CP-element group 283: 	 branch_block_stmt_655/if_stmt_2096_else_link/$entry
      -- 
    ca_5394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2081_inst_ack_1, ack => zeropad3D_CP_2067_elements(283)); -- 
    branch_req_5402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(283), ack => if_stmt_2096_branch_req_0); -- 
    -- CP-element group 284:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	938 
    -- CP-element group 284: 	939 
    -- CP-element group 284: 	941 
    -- CP-element group 284: 	942 
    -- CP-element group 284: 	944 
    -- CP-element group 284: 	945 
    -- CP-element group 284:  members (40) 
      -- CP-element group 284: 	 branch_block_stmt_655/merge_stmt_2102__exit__
      -- CP-element group 284: 	 branch_block_stmt_655/assign_stmt_2108__entry__
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607
      -- CP-element group 284: 	 branch_block_stmt_655/assign_stmt_2108__exit__
      -- CP-element group 284: 	 branch_block_stmt_655/if_stmt_2096_if_link/$exit
      -- CP-element group 284: 	 branch_block_stmt_655/if_stmt_2096_if_link/if_choice_transition
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xend555_ifx_xthen565
      -- CP-element group 284: 	 branch_block_stmt_655/assign_stmt_2108/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/assign_stmt_2108/$exit
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xend555_ifx_xthen565_PhiReq/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xend555_ifx_xthen565_PhiReq/$exit
      -- CP-element group 284: 	 branch_block_stmt_655/merge_stmt_2102_PhiReqMerge
      -- CP-element group 284: 	 branch_block_stmt_655/merge_stmt_2102_PhiAck/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/merge_stmt_2102_PhiAck/$exit
      -- CP-element group 284: 	 branch_block_stmt_655/merge_stmt_2102_PhiAck/dummy
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/Update/cr
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/Update/cr
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2096_branch_ack_1, ack => zeropad3D_CP_2067_elements(284)); -- 
    rr_11759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(284), ack => type_cast_2199_inst_req_0); -- 
    cr_11764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(284), ack => type_cast_2199_inst_req_1); -- 
    rr_11782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(284), ack => type_cast_2208_inst_req_0); -- 
    cr_11787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(284), ack => type_cast_2208_inst_req_1); -- 
    rr_11805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(284), ack => type_cast_2214_inst_req_0); -- 
    cr_11810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(284), ack => type_cast_2214_inst_req_1); -- 
    -- CP-element group 285:  fork  transition  place  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285: 	287 
    -- CP-element group 285: 	288 
    -- CP-element group 285: 	289 
    -- CP-element group 285: 	291 
    -- CP-element group 285: 	294 
    -- CP-element group 285: 	296 
    -- CP-element group 285: 	297 
    -- CP-element group 285: 	298 
    -- CP-element group 285: 	300 
    -- CP-element group 285:  members (54) 
      -- CP-element group 285: 	 branch_block_stmt_655/merge_stmt_2110__exit__
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188__entry__
      -- CP-element group 285: 	 branch_block_stmt_655/if_stmt_2096_else_link/$exit
      -- CP-element group 285: 	 branch_block_stmt_655/if_stmt_2096_else_link/else_choice_transition
      -- CP-element group 285: 	 branch_block_stmt_655/ifx_xend555_ifx_xelse570
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_sample_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_update_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_Sample/rr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_Update/cr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_sample_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_update_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_word_address_calculated
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_root_address_calculated
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Sample/word_access_start/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Sample/word_access_start/word_0/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Sample/word_access_start/word_0/rr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/word_access_complete/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/word_access_complete/word_0/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/word_access_complete/word_0/cr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_update_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_Update/cr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_update_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_Update/cr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_update_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_Update/cr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_sample_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_update_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_word_address_calculated
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_root_address_calculated
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Sample/word_access_start/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Sample/word_access_start/word_0/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Sample/word_access_start/word_0/rr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/word_access_complete/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/word_access_complete/word_0/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/word_access_complete/word_0/cr
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_update_start_
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_Update/cr
      -- CP-element group 285: 	 branch_block_stmt_655/ifx_xend555_ifx_xelse570_PhiReq/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/ifx_xend555_ifx_xelse570_PhiReq/$exit
      -- CP-element group 285: 	 branch_block_stmt_655/merge_stmt_2110_PhiReqMerge
      -- CP-element group 285: 	 branch_block_stmt_655/merge_stmt_2110_PhiAck/$entry
      -- CP-element group 285: 	 branch_block_stmt_655/merge_stmt_2110_PhiAck/$exit
      -- CP-element group 285: 	 branch_block_stmt_655/merge_stmt_2110_PhiAck/dummy
      -- 
    else_choice_transition_5411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2096_branch_ack_0, ack => zeropad3D_CP_2067_elements(285)); -- 
    rr_5427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => type_cast_2120_inst_req_0); -- 
    cr_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => type_cast_2120_inst_req_1); -- 
    rr_5449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => LOAD_col_high_2123_load_0_req_0); -- 
    cr_5460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => LOAD_col_high_2123_load_0_req_1); -- 
    cr_5479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => type_cast_2127_inst_req_1); -- 
    cr_5493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => type_cast_2147_inst_req_1); -- 
    cr_5507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => type_cast_2164_inst_req_1); -- 
    rr_5524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => LOAD_row_high_2167_load_0_req_0); -- 
    cr_5535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => LOAD_row_high_2167_load_0_req_1); -- 
    cr_5554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(285), ack => type_cast_2171_inst_req_1); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_Sample/ra
      -- 
    ra_5428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2120_inst_ack_0, ack => zeropad3D_CP_2067_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	292 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2120_Update/ca
      -- 
    ca_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2120_inst_ack_1, ack => zeropad3D_CP_2067_elements(287)); -- 
    -- CP-element group 288:  transition  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: successors 
    -- CP-element group 288:  members (5) 
      -- CP-element group 288: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Sample/word_access_start/$exit
      -- CP-element group 288: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Sample/word_access_start/word_0/$exit
      -- CP-element group 288: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Sample/word_access_start/word_0/ra
      -- 
    ra_5450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2123_load_0_ack_0, ack => zeropad3D_CP_2067_elements(288)); -- 
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	285 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (12) 
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/word_access_complete/$exit
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/word_access_complete/word_0/$exit
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/word_access_complete/word_0/ca
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/LOAD_col_high_2123_Merge/$entry
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/LOAD_col_high_2123_Merge/$exit
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/LOAD_col_high_2123_Merge/merge_req
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_col_high_2123_Update/LOAD_col_high_2123_Merge/merge_ack
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_Sample/rr
      -- 
    ca_5461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2123_load_0_ack_1, ack => zeropad3D_CP_2067_elements(289)); -- 
    rr_5474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(289), ack => type_cast_2127_inst_req_0); -- 
    -- CP-element group 290:  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_Sample/ra
      -- 
    ra_5475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2127_inst_ack_0, ack => zeropad3D_CP_2067_elements(290)); -- 
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	285 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_Update/$exit
      -- CP-element group 291: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2127_Update/ca
      -- 
    ca_5480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2127_inst_ack_1, ack => zeropad3D_CP_2067_elements(291)); -- 
    -- CP-element group 292:  join  transition  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	287 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_Sample/rr
      -- 
    rr_5488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(292), ack => type_cast_2147_inst_req_0); -- 
    zeropad3D_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(287) & zeropad3D_CP_2067_elements(291);
      gj_zeropad3D_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_Sample/ra
      -- 
    ra_5489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_0, ack => zeropad3D_CP_2067_elements(293)); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	285 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2147_Update/ca
      -- CP-element group 294: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_Sample/rr
      -- 
    ca_5494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2147_inst_ack_1, ack => zeropad3D_CP_2067_elements(294)); -- 
    rr_5502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(294), ack => type_cast_2164_inst_req_0); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_Sample/ra
      -- 
    ra_5503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2164_inst_ack_0, ack => zeropad3D_CP_2067_elements(295)); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	285 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	301 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2164_Update/ca
      -- 
    ca_5508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2164_inst_ack_1, ack => zeropad3D_CP_2067_elements(296)); -- 
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	285 
    -- CP-element group 297: successors 
    -- CP-element group 297:  members (5) 
      -- CP-element group 297: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Sample/word_access_start/$exit
      -- CP-element group 297: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Sample/word_access_start/word_0/$exit
      -- CP-element group 297: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Sample/word_access_start/word_0/ra
      -- 
    ra_5525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2167_load_0_ack_0, ack => zeropad3D_CP_2067_elements(297)); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	285 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (12) 
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/word_access_complete/$exit
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/word_access_complete/word_0/$exit
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/word_access_complete/word_0/ca
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/LOAD_row_high_2167_Merge/$entry
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/LOAD_row_high_2167_Merge/$exit
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/LOAD_row_high_2167_Merge/merge_req
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/LOAD_row_high_2167_Update/LOAD_row_high_2167_Merge/merge_ack
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_Sample/rr
      -- 
    ca_5536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2167_load_0_ack_1, ack => zeropad3D_CP_2067_elements(298)); -- 
    rr_5549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(298), ack => type_cast_2171_inst_req_0); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_Sample/ra
      -- 
    ra_5550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2171_inst_ack_0, ack => zeropad3D_CP_2067_elements(299)); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	285 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/type_cast_2171_Update/ca
      -- 
    ca_5555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2171_inst_ack_1, ack => zeropad3D_CP_2067_elements(300)); -- 
    -- CP-element group 301:  branch  join  transition  place  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	296 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (10) 
      -- CP-element group 301: 	 branch_block_stmt_655/if_stmt_2189__entry__
      -- CP-element group 301: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188__exit__
      -- CP-element group 301: 	 branch_block_stmt_655/assign_stmt_2116_to_assign_stmt_2188/$exit
      -- CP-element group 301: 	 branch_block_stmt_655/if_stmt_2189_dead_link/$entry
      -- CP-element group 301: 	 branch_block_stmt_655/if_stmt_2189_eval_test/$entry
      -- CP-element group 301: 	 branch_block_stmt_655/if_stmt_2189_eval_test/$exit
      -- CP-element group 301: 	 branch_block_stmt_655/if_stmt_2189_eval_test/branch_req
      -- CP-element group 301: 	 branch_block_stmt_655/R_cmp598_2190_place
      -- CP-element group 301: 	 branch_block_stmt_655/if_stmt_2189_if_link/$entry
      -- CP-element group 301: 	 branch_block_stmt_655/if_stmt_2189_else_link/$entry
      -- 
    branch_req_5563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(301), ack => if_stmt_2189_branch_req_0); -- 
    zeropad3D_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(296) & zeropad3D_CP_2067_elements(300);
      gj_zeropad3D_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  fork  transition  place  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	953 
    -- CP-element group 302: 	954 
    -- CP-element group 302: 	956 
    -- CP-element group 302: 	957 
    -- CP-element group 302: 	959 
    -- CP-element group 302: 	960 
    -- CP-element group 302:  members (28) 
      -- CP-element group 302: 	 branch_block_stmt_655/if_stmt_2189_if_link/$exit
      -- CP-element group 302: 	 branch_block_stmt_655/if_stmt_2189_if_link/if_choice_transition
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/Sample/rr
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/Update/cr
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/Sample/rr
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/Update/cr
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/Sample/rr
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2189_branch_ack_1, ack => zeropad3D_CP_2067_elements(302)); -- 
    rr_11838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(302), ack => type_cast_2221_inst_req_0); -- 
    cr_11843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(302), ack => type_cast_2221_inst_req_1); -- 
    rr_11861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(302), ack => type_cast_2225_inst_req_0); -- 
    cr_11866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(302), ack => type_cast_2225_inst_req_1); -- 
    rr_11884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(302), ack => type_cast_2229_inst_req_0); -- 
    cr_11889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(302), ack => type_cast_2229_inst_req_1); -- 
    -- CP-element group 303:  fork  transition  place  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	930 
    -- CP-element group 303: 	931 
    -- CP-element group 303: 	932 
    -- CP-element group 303: 	934 
    -- CP-element group 303: 	935 
    -- CP-element group 303:  members (22) 
      -- CP-element group 303: 	 branch_block_stmt_655/if_stmt_2189_else_link/$exit
      -- CP-element group 303: 	 branch_block_stmt_655/if_stmt_2189_else_link/else_choice_transition
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2196/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/Update/cr
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/Sample/rr
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2189_branch_ack_0, ack => zeropad3D_CP_2067_elements(303)); -- 
    rr_11710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(303), ack => type_cast_2206_inst_req_0); -- 
    cr_11715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(303), ack => type_cast_2206_inst_req_1); -- 
    rr_11733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(303), ack => type_cast_2212_inst_req_0); -- 
    cr_11738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(303), ack => type_cast_2212_inst_req_1); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	966 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_sample_completed_
      -- CP-element group 304: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_Sample/$exit
      -- CP-element group 304: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_Sample/ra
      -- 
    ra_5586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2233_inst_ack_0, ack => zeropad3D_CP_2067_elements(304)); -- 
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	966 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	326 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_update_completed_
      -- CP-element group 305: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_Update/$exit
      -- CP-element group 305: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_Update/ca
      -- 
    ca_5591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2233_inst_ack_1, ack => zeropad3D_CP_2067_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	966 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_Sample/ra
      -- 
    ra_5600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2243_inst_ack_0, ack => zeropad3D_CP_2067_elements(306)); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	966 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	326 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_update_completed_
      -- CP-element group 307: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_Update/ca
      -- 
    ca_5605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2243_inst_ack_1, ack => zeropad3D_CP_2067_elements(307)); -- 
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	966 
    -- CP-element group 308: successors 
    -- CP-element group 308:  members (5) 
      -- CP-element group 308: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_sample_completed_
      -- CP-element group 308: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Sample/$exit
      -- CP-element group 308: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Sample/word_access_start/$exit
      -- CP-element group 308: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Sample/word_access_start/word_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Sample/word_access_start/word_0/ra
      -- 
    ra_5622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2252_load_0_ack_0, ack => zeropad3D_CP_2067_elements(308)); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	966 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	322 
    -- CP-element group 309:  members (12) 
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_Sample/rr
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_update_completed_
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/$exit
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/word_access_complete/$exit
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/word_access_complete/word_0/$exit
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/word_access_complete/word_0/ca
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/LOAD_pad_2252_Merge/$entry
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/LOAD_pad_2252_Merge/$exit
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/LOAD_pad_2252_Merge/merge_req
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/LOAD_pad_2252_Merge/merge_ack
      -- CP-element group 309: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_sample_start_
      -- 
    ca_5633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2252_load_0_ack_1, ack => zeropad3D_CP_2067_elements(309)); -- 
    rr_5787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(309), ack => type_cast_2282_inst_req_0); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	966 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (5) 
      -- CP-element group 310: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Sample/word_access_start/$exit
      -- CP-element group 310: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Sample/word_access_start/word_0/$exit
      -- CP-element group 310: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Sample/word_access_start/word_0/ra
      -- 
    ra_5655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_2255_load_0_ack_0, ack => zeropad3D_CP_2067_elements(310)); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	966 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	316 
    -- CP-element group 311:  members (12) 
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/word_access_complete/$exit
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/word_access_complete/word_0/$exit
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/word_access_complete/word_0/ca
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/LOAD_depth_high_2255_Merge/$entry
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/LOAD_depth_high_2255_Merge/$exit
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/LOAD_depth_high_2255_Merge/merge_req
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/LOAD_depth_high_2255_Merge/merge_ack
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_sample_start_
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_Sample/rr
      -- 
    ca_5666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_2255_load_0_ack_1, ack => zeropad3D_CP_2067_elements(311)); -- 
    rr_5745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(311), ack => type_cast_2265_inst_req_0); -- 
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	966 
    -- CP-element group 312: successors 
    -- CP-element group 312:  members (5) 
      -- CP-element group 312: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Sample/word_access_start/$exit
      -- CP-element group 312: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Sample/word_access_start/word_0/$exit
      -- CP-element group 312: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Sample/word_access_start/word_0/ra
      -- 
    ra_5688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_2258_load_0_ack_0, ack => zeropad3D_CP_2067_elements(312)); -- 
    -- CP-element group 313:  fork  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	966 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	318 
    -- CP-element group 313: 	324 
    -- CP-element group 313:  members (15) 
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_Sample/rr
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/word_access_complete/$exit
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/word_access_complete/word_0/$exit
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/word_access_complete/word_0/ca
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/LOAD_out_depth_high_2258_Merge/$entry
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/LOAD_out_depth_high_2258_Merge/$exit
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/LOAD_out_depth_high_2258_Merge/merge_req
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/LOAD_out_depth_high_2258_Merge/merge_ack
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_Sample/rr
      -- 
    ca_5699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_2258_load_0_ack_1, ack => zeropad3D_CP_2067_elements(313)); -- 
    rr_5759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(313), ack => type_cast_2269_inst_req_0); -- 
    rr_5801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(313), ack => type_cast_2286_inst_req_0); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	966 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (5) 
      -- CP-element group 314: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_sample_completed_
      -- CP-element group 314: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Sample/word_access_start/$exit
      -- CP-element group 314: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Sample/word_access_start/word_0/$exit
      -- CP-element group 314: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Sample/word_access_start/word_0/ra
      -- 
    ra_5721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_2261_load_0_ack_0, ack => zeropad3D_CP_2067_elements(314)); -- 
    -- CP-element group 315:  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	966 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	320 
    -- CP-element group 315:  members (12) 
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_update_completed_
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/$exit
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/word_access_complete/$exit
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/word_access_complete/word_0/$exit
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/word_access_complete/word_0/ca
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/LOAD_out_col_high_2261_Merge/$entry
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/LOAD_out_col_high_2261_Merge/$exit
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/LOAD_out_col_high_2261_Merge/merge_req
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/LOAD_out_col_high_2261_Merge/merge_ack
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_sample_start_
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_Sample/$entry
      -- CP-element group 315: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_Sample/rr
      -- 
    ca_5732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_2261_load_0_ack_1, ack => zeropad3D_CP_2067_elements(315)); -- 
    rr_5773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(315), ack => type_cast_2273_inst_req_0); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	311 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_sample_completed_
      -- CP-element group 316: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_Sample/ra
      -- 
    ra_5746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2265_inst_ack_0, ack => zeropad3D_CP_2067_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	966 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	326 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_update_completed_
      -- CP-element group 317: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_Update/$exit
      -- CP-element group 317: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_Update/ca
      -- 
    ca_5751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2265_inst_ack_1, ack => zeropad3D_CP_2067_elements(317)); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	313 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_Sample/ra
      -- 
    ra_5760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2269_inst_ack_0, ack => zeropad3D_CP_2067_elements(318)); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	966 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	326 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_Update/ca
      -- 
    ca_5765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2269_inst_ack_1, ack => zeropad3D_CP_2067_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	315 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_Sample/ra
      -- 
    ra_5774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2273_inst_ack_0, ack => zeropad3D_CP_2067_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	966 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	326 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_Update/ca
      -- 
    ca_5779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2273_inst_ack_1, ack => zeropad3D_CP_2067_elements(321)); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	309 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_Sample/ra
      -- CP-element group 322: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_Sample/$exit
      -- CP-element group 322: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_sample_completed_
      -- 
    ra_5788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2282_inst_ack_0, ack => zeropad3D_CP_2067_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	966 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	326 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_Update/$exit
      -- CP-element group 323: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_Update/ca
      -- CP-element group 323: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_update_completed_
      -- 
    ca_5793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2282_inst_ack_1, ack => zeropad3D_CP_2067_elements(323)); -- 
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	313 
    -- CP-element group 324: successors 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_Sample/ra
      -- 
    ra_5802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2286_inst_ack_0, ack => zeropad3D_CP_2067_elements(324)); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	966 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_Update/ca
      -- CP-element group 325: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_Update/$exit
      -- 
    ca_5807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2286_inst_ack_1, ack => zeropad3D_CP_2067_elements(325)); -- 
    -- CP-element group 326:  join  fork  transition  place  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	305 
    -- CP-element group 326: 	307 
    -- CP-element group 326: 	317 
    -- CP-element group 326: 	319 
    -- CP-element group 326: 	321 
    -- CP-element group 326: 	323 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	977 
    -- CP-element group 326: 	978 
    -- CP-element group 326: 	979 
    -- CP-element group 326: 	981 
    -- CP-element group 326: 	982 
    -- CP-element group 326:  members (22) 
      -- CP-element group 326: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328__exit__
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672
      -- CP-element group 326: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/$exit
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2331/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/Update/cr
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/Update/cr
      -- 
    rr_11997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(326), ack => type_cast_2341_inst_req_0); -- 
    cr_12002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(326), ack => type_cast_2341_inst_req_1); -- 
    rr_12020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(326), ack => type_cast_2347_inst_req_0); -- 
    cr_12025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(326), ack => type_cast_2347_inst_req_1); -- 
    zeropad3D_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(305) & zeropad3D_CP_2067_elements(307) & zeropad3D_CP_2067_elements(317) & zeropad3D_CP_2067_elements(319) & zeropad3D_CP_2067_elements(321) & zeropad3D_CP_2067_elements(323) & zeropad3D_CP_2067_elements(325);
      gj_zeropad3D_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	989 
    -- CP-element group 327: successors 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_Sample/ra
      -- CP-element group 327: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_Sample/$exit
      -- 
    ra_5819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2354_inst_ack_0, ack => zeropad3D_CP_2067_elements(327)); -- 
    -- CP-element group 328:  branch  transition  place  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	989 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328: 	330 
    -- CP-element group 328:  members (13) 
      -- CP-element group 328: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362__exit__
      -- CP-element group 328: 	 branch_block_stmt_655/if_stmt_2363__entry__
      -- CP-element group 328: 	 branch_block_stmt_655/if_stmt_2363_dead_link/$entry
      -- CP-element group 328: 	 branch_block_stmt_655/if_stmt_2363_eval_test/$entry
      -- CP-element group 328: 	 branch_block_stmt_655/if_stmt_2363_eval_test/$exit
      -- CP-element group 328: 	 branch_block_stmt_655/if_stmt_2363_eval_test/branch_req
      -- CP-element group 328: 	 branch_block_stmt_655/if_stmt_2363_if_link/$entry
      -- CP-element group 328: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_655/if_stmt_2363_else_link/$entry
      -- CP-element group 328: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_Update/ca
      -- CP-element group 328: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/$exit
      -- CP-element group 328: 	 branch_block_stmt_655/R_cmp677_2364_place
      -- CP-element group 328: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_Update/$exit
      -- 
    ca_5824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2354_inst_ack_1, ack => zeropad3D_CP_2067_elements(328)); -- 
    branch_req_5832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(328), ack => if_stmt_2363_branch_req_0); -- 
    -- CP-element group 329:  transition  place  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	990 
    -- CP-element group 329:  members (5) 
      -- CP-element group 329: 	 branch_block_stmt_655/whilex_xbody672_ifx_xthen707
      -- CP-element group 329: 	 branch_block_stmt_655/if_stmt_2363_if_link/$exit
      -- CP-element group 329: 	 branch_block_stmt_655/if_stmt_2363_if_link/if_choice_transition
      -- CP-element group 329: 	 branch_block_stmt_655/whilex_xbody672_ifx_xthen707_PhiReq/$entry
      -- CP-element group 329: 	 branch_block_stmt_655/whilex_xbody672_ifx_xthen707_PhiReq/$exit
      -- 
    if_choice_transition_5837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2363_branch_ack_1, ack => zeropad3D_CP_2067_elements(329)); -- 
    -- CP-element group 330:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	328 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330: 	332 
    -- CP-element group 330: 	334 
    -- CP-element group 330:  members (27) 
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394__entry__
      -- CP-element group 330: 	 branch_block_stmt_655/merge_stmt_2369__exit__
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_update_start_
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_update_start_
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_Update/cr
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_word_address_calculated
      -- CP-element group 330: 	 branch_block_stmt_655/whilex_xbody672_lorx_xlhsx_xfalse679
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_root_address_calculated
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Sample/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/if_stmt_2363_else_link/$exit
      -- CP-element group 330: 	 branch_block_stmt_655/if_stmt_2363_else_link/else_choice_transition
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_sample_start_
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/word_access_complete/word_0/cr
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/word_access_complete/word_0/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/word_access_complete/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Sample/word_access_start/word_0/rr
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Sample/word_access_start/word_0/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Sample/word_access_start/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/whilex_xbody672_lorx_xlhsx_xfalse679_PhiReq/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/whilex_xbody672_lorx_xlhsx_xfalse679_PhiReq/$exit
      -- CP-element group 330: 	 branch_block_stmt_655/merge_stmt_2369_PhiReqMerge
      -- CP-element group 330: 	 branch_block_stmt_655/merge_stmt_2369_PhiAck/$entry
      -- CP-element group 330: 	 branch_block_stmt_655/merge_stmt_2369_PhiAck/$exit
      -- CP-element group 330: 	 branch_block_stmt_655/merge_stmt_2369_PhiAck/dummy
      -- 
    else_choice_transition_5841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2363_branch_ack_0, ack => zeropad3D_CP_2067_elements(330)); -- 
    cr_5892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(330), ack => type_cast_2375_inst_req_1); -- 
    cr_5873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(330), ack => LOAD_row_high_2371_load_0_req_1); -- 
    rr_5862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(330), ack => LOAD_row_high_2371_load_0_req_0); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331:  members (5) 
      -- CP-element group 331: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Sample/word_access_start/word_0/ra
      -- CP-element group 331: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Sample/word_access_start/word_0/$exit
      -- CP-element group 331: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Sample/word_access_start/$exit
      -- CP-element group 331: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Sample/$exit
      -- 
    ra_5863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2371_load_0_ack_0, ack => zeropad3D_CP_2067_elements(331)); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (12) 
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/LOAD_row_high_2371_Merge/merge_ack
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_Sample/rr
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/LOAD_row_high_2371_Merge/merge_req
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/LOAD_row_high_2371_Merge/$exit
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/LOAD_row_high_2371_Merge/$entry
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/word_access_complete/word_0/ca
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/word_access_complete/word_0/$exit
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/word_access_complete/$exit
      -- CP-element group 332: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/LOAD_row_high_2371_Update/$exit
      -- 
    ca_5874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2371_load_0_ack_1, ack => zeropad3D_CP_2067_elements(332)); -- 
    rr_5887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(332), ack => type_cast_2375_inst_req_0); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_Sample/ra
      -- 
    ra_5888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2375_inst_ack_0, ack => zeropad3D_CP_2067_elements(333)); -- 
    -- CP-element group 334:  branch  transition  place  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	330 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (13) 
      -- CP-element group 334: 	 branch_block_stmt_655/if_stmt_2395__entry__
      -- CP-element group 334: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394__exit__
      -- CP-element group 334: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/type_cast_2375_Update/ca
      -- CP-element group 334: 	 branch_block_stmt_655/if_stmt_2395_dead_link/$entry
      -- CP-element group 334: 	 branch_block_stmt_655/if_stmt_2395_eval_test/$entry
      -- CP-element group 334: 	 branch_block_stmt_655/if_stmt_2395_eval_test/$exit
      -- CP-element group 334: 	 branch_block_stmt_655/if_stmt_2395_eval_test/branch_req
      -- CP-element group 334: 	 branch_block_stmt_655/if_stmt_2395_if_link/$entry
      -- CP-element group 334: 	 branch_block_stmt_655/if_stmt_2395_else_link/$entry
      -- CP-element group 334: 	 branch_block_stmt_655/R_cmp688_2396_place
      -- CP-element group 334: 	 branch_block_stmt_655/assign_stmt_2372_to_assign_stmt_2394/$exit
      -- 
    ca_5893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2375_inst_ack_1, ack => zeropad3D_CP_2067_elements(334)); -- 
    branch_req_5901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(334), ack => if_stmt_2395_branch_req_0); -- 
    -- CP-element group 335:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: 	338 
    -- CP-element group 335:  members (18) 
      -- CP-element group 335: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413__entry__
      -- CP-element group 335: 	 branch_block_stmt_655/merge_stmt_2401__exit__
      -- CP-element group 335: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_update_start_
      -- CP-element group 335: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_655/if_stmt_2395_if_link/$exit
      -- CP-element group 335: 	 branch_block_stmt_655/if_stmt_2395_if_link/if_choice_transition
      -- CP-element group 335: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/$entry
      -- CP-element group 335: 	 branch_block_stmt_655/lorx_xlhsx_xfalse679_lorx_xlhsx_xfalse690
      -- CP-element group 335: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_655/lorx_xlhsx_xfalse679_lorx_xlhsx_xfalse690_PhiReq/$entry
      -- CP-element group 335: 	 branch_block_stmt_655/lorx_xlhsx_xfalse679_lorx_xlhsx_xfalse690_PhiReq/$exit
      -- CP-element group 335: 	 branch_block_stmt_655/merge_stmt_2401_PhiReqMerge
      -- CP-element group 335: 	 branch_block_stmt_655/merge_stmt_2401_PhiAck/$entry
      -- CP-element group 335: 	 branch_block_stmt_655/merge_stmt_2401_PhiAck/$exit
      -- CP-element group 335: 	 branch_block_stmt_655/merge_stmt_2401_PhiAck/dummy
      -- 
    if_choice_transition_5906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2395_branch_ack_1, ack => zeropad3D_CP_2067_elements(335)); -- 
    rr_5923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(335), ack => type_cast_2405_inst_req_0); -- 
    cr_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(335), ack => type_cast_2405_inst_req_1); -- 
    -- CP-element group 336:  transition  place  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	990 
    -- CP-element group 336:  members (5) 
      -- CP-element group 336: 	 branch_block_stmt_655/if_stmt_2395_else_link/$exit
      -- CP-element group 336: 	 branch_block_stmt_655/if_stmt_2395_else_link/else_choice_transition
      -- CP-element group 336: 	 branch_block_stmt_655/lorx_xlhsx_xfalse679_ifx_xthen707
      -- CP-element group 336: 	 branch_block_stmt_655/lorx_xlhsx_xfalse679_ifx_xthen707_PhiReq/$entry
      -- CP-element group 336: 	 branch_block_stmt_655/lorx_xlhsx_xfalse679_ifx_xthen707_PhiReq/$exit
      -- 
    else_choice_transition_5910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2395_branch_ack_0, ack => zeropad3D_CP_2067_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_Sample/ra
      -- CP-element group 337: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_sample_completed_
      -- 
    ra_5924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2405_inst_ack_0, ack => zeropad3D_CP_2067_elements(337)); -- 
    -- CP-element group 338:  branch  transition  place  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	335 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (13) 
      -- CP-element group 338: 	 branch_block_stmt_655/if_stmt_2414__entry__
      -- CP-element group 338: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413__exit__
      -- CP-element group 338: 	 branch_block_stmt_655/R_cmp695_2415_place
      -- CP-element group 338: 	 branch_block_stmt_655/if_stmt_2414_if_link/$entry
      -- CP-element group 338: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_655/if_stmt_2414_else_link/$entry
      -- CP-element group 338: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/$exit
      -- CP-element group 338: 	 branch_block_stmt_655/if_stmt_2414_eval_test/branch_req
      -- CP-element group 338: 	 branch_block_stmt_655/if_stmt_2414_eval_test/$exit
      -- CP-element group 338: 	 branch_block_stmt_655/if_stmt_2414_eval_test/$entry
      -- CP-element group 338: 	 branch_block_stmt_655/if_stmt_2414_dead_link/$entry
      -- CP-element group 338: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_Update/ca
      -- CP-element group 338: 	 branch_block_stmt_655/assign_stmt_2406_to_assign_stmt_2413/type_cast_2405_Update/$exit
      -- 
    ca_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2405_inst_ack_1, ack => zeropad3D_CP_2067_elements(338)); -- 
    branch_req_5937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(338), ack => if_stmt_2414_branch_req_0); -- 
    -- CP-element group 339:  transition  place  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	990 
    -- CP-element group 339:  members (5) 
      -- CP-element group 339: 	 branch_block_stmt_655/if_stmt_2414_if_link/$exit
      -- CP-element group 339: 	 branch_block_stmt_655/if_stmt_2414_if_link/if_choice_transition
      -- CP-element group 339: 	 branch_block_stmt_655/lorx_xlhsx_xfalse690_ifx_xthen707
      -- CP-element group 339: 	 branch_block_stmt_655/lorx_xlhsx_xfalse690_ifx_xthen707_PhiReq/$entry
      -- CP-element group 339: 	 branch_block_stmt_655/lorx_xlhsx_xfalse690_ifx_xthen707_PhiReq/$exit
      -- 
    if_choice_transition_5942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2414_branch_ack_1, ack => zeropad3D_CP_2067_elements(339)); -- 
    -- CP-element group 340:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340: 	342 
    -- CP-element group 340: 	344 
    -- CP-element group 340:  members (27) 
      -- CP-element group 340: 	 branch_block_stmt_655/merge_stmt_2420__exit__
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439__entry__
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_word_address_calculated
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_root_address_calculated
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_Update/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/if_stmt_2414_else_link/$exit
      -- CP-element group 340: 	 branch_block_stmt_655/if_stmt_2414_else_link/else_choice_transition
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_Update/cr
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Sample/word_access_start/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/lorx_xlhsx_xfalse690_lorx_xlhsx_xfalse697
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Sample/word_access_start/word_0/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/word_access_complete/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Sample/word_access_start/word_0/rr
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_update_start_
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/word_access_complete/word_0/cr
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_update_start_
      -- CP-element group 340: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/word_access_complete/word_0/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/lorx_xlhsx_xfalse690_lorx_xlhsx_xfalse697_PhiReq/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/lorx_xlhsx_xfalse690_lorx_xlhsx_xfalse697_PhiReq/$exit
      -- CP-element group 340: 	 branch_block_stmt_655/merge_stmt_2420_PhiReqMerge
      -- CP-element group 340: 	 branch_block_stmt_655/merge_stmt_2420_PhiAck/$entry
      -- CP-element group 340: 	 branch_block_stmt_655/merge_stmt_2420_PhiAck/$exit
      -- CP-element group 340: 	 branch_block_stmt_655/merge_stmt_2420_PhiAck/dummy
      -- 
    else_choice_transition_5946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2414_branch_ack_0, ack => zeropad3D_CP_2067_elements(340)); -- 
    cr_5997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(340), ack => type_cast_2426_inst_req_1); -- 
    rr_5967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(340), ack => LOAD_col_high_2422_load_0_req_0); -- 
    cr_5978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(340), ack => LOAD_col_high_2422_load_0_req_1); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341:  members (5) 
      -- CP-element group 341: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Sample/word_access_start/word_0/$exit
      -- CP-element group 341: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Sample/word_access_start/$exit
      -- CP-element group 341: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Sample/word_access_start/word_0/ra
      -- 
    ra_5968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2422_load_0_ack_0, ack => zeropad3D_CP_2067_elements(341)); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (12) 
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/LOAD_col_high_2422_Merge/$entry
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/LOAD_col_high_2422_Merge/$exit
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/LOAD_col_high_2422_Merge/merge_req
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_Sample/rr
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/LOAD_col_high_2422_Merge/merge_ack
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/word_access_complete/$exit
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/word_access_complete/word_0/ca
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/LOAD_col_high_2422_Update/word_access_complete/word_0/$exit
      -- CP-element group 342: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_sample_start_
      -- 
    ca_5979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2422_load_0_ack_1, ack => zeropad3D_CP_2067_elements(342)); -- 
    rr_5992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(342), ack => type_cast_2426_inst_req_0); -- 
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_Sample/ra
      -- CP-element group 343: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_sample_completed_
      -- 
    ra_5993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2426_inst_ack_0, ack => zeropad3D_CP_2067_elements(343)); -- 
    -- CP-element group 344:  branch  transition  place  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	340 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (13) 
      -- CP-element group 344: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439__exit__
      -- CP-element group 344: 	 branch_block_stmt_655/if_stmt_2440__entry__
      -- CP-element group 344: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_Update/ca
      -- CP-element group 344: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/$exit
      -- CP-element group 344: 	 branch_block_stmt_655/assign_stmt_2423_to_assign_stmt_2439/type_cast_2426_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_655/if_stmt_2440_dead_link/$entry
      -- CP-element group 344: 	 branch_block_stmt_655/if_stmt_2440_eval_test/$entry
      -- CP-element group 344: 	 branch_block_stmt_655/if_stmt_2440_eval_test/$exit
      -- CP-element group 344: 	 branch_block_stmt_655/if_stmt_2440_eval_test/branch_req
      -- CP-element group 344: 	 branch_block_stmt_655/R_cmp705_2441_place
      -- CP-element group 344: 	 branch_block_stmt_655/if_stmt_2440_if_link/$entry
      -- CP-element group 344: 	 branch_block_stmt_655/if_stmt_2440_else_link/$entry
      -- 
    ca_5998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2426_inst_ack_1, ack => zeropad3D_CP_2067_elements(344)); -- 
    branch_req_6006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(344), ack => if_stmt_2440_branch_req_0); -- 
    -- CP-element group 345:  fork  transition  place  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	361 
    -- CP-element group 345: 	362 
    -- CP-element group 345: 	364 
    -- CP-element group 345: 	366 
    -- CP-element group 345: 	368 
    -- CP-element group 345: 	370 
    -- CP-element group 345: 	372 
    -- CP-element group 345: 	374 
    -- CP-element group 345: 	376 
    -- CP-element group 345: 	379 
    -- CP-element group 345:  members (46) 
      -- CP-element group 345: 	 branch_block_stmt_655/merge_stmt_2504__exit__
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609__entry__
      -- CP-element group 345: 	 branch_block_stmt_655/if_stmt_2440_if_link/$exit
      -- CP-element group 345: 	 branch_block_stmt_655/if_stmt_2440_if_link/if_choice_transition
      -- CP-element group 345: 	 branch_block_stmt_655/lorx_xlhsx_xfalse697_ifx_xelse728
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_sample_start_
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_update_start_
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_Sample/rr
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_Update/cr
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_update_start_
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_Update/cr
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_update_start_
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_update_start
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_Update/req
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_complete/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_complete/req
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_update_start_
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/word_access_complete/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/word_access_complete/word_0/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/word_access_complete/word_0/cr
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_update_start_
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_Update/cr
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_update_start_
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_update_start
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_Update/req
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_complete/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_complete/req
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_update_start_
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Update/word_access_complete/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Update/word_access_complete/word_0/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Update/word_access_complete/word_0/cr
      -- CP-element group 345: 	 branch_block_stmt_655/lorx_xlhsx_xfalse697_ifx_xelse728_PhiReq/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/lorx_xlhsx_xfalse697_ifx_xelse728_PhiReq/$exit
      -- CP-element group 345: 	 branch_block_stmt_655/merge_stmt_2504_PhiReqMerge
      -- CP-element group 345: 	 branch_block_stmt_655/merge_stmt_2504_PhiAck/$entry
      -- CP-element group 345: 	 branch_block_stmt_655/merge_stmt_2504_PhiAck/$exit
      -- CP-element group 345: 	 branch_block_stmt_655/merge_stmt_2504_PhiAck/dummy
      -- 
    if_choice_transition_6011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2440_branch_ack_1, ack => zeropad3D_CP_2067_elements(345)); -- 
    rr_6169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => type_cast_2508_inst_req_0); -- 
    cr_6174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => type_cast_2508_inst_req_1); -- 
    cr_6188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => type_cast_2572_inst_req_1); -- 
    req_6219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => array_obj_ref_2578_index_offset_req_1); -- 
    req_6234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => addr_of_2579_final_reg_req_1); -- 
    cr_6279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => ptr_deref_2583_load_0_req_1); -- 
    cr_6298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => type_cast_2597_inst_req_1); -- 
    req_6329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => array_obj_ref_2603_index_offset_req_1); -- 
    req_6344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => addr_of_2604_final_reg_req_1); -- 
    cr_6394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(345), ack => ptr_deref_2607_store_0_req_1); -- 
    -- CP-element group 346:  transition  place  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	990 
    -- CP-element group 346:  members (5) 
      -- CP-element group 346: 	 branch_block_stmt_655/if_stmt_2440_else_link/$exit
      -- CP-element group 346: 	 branch_block_stmt_655/if_stmt_2440_else_link/else_choice_transition
      -- CP-element group 346: 	 branch_block_stmt_655/lorx_xlhsx_xfalse697_ifx_xthen707
      -- CP-element group 346: 	 branch_block_stmt_655/lorx_xlhsx_xfalse697_ifx_xthen707_PhiReq/$entry
      -- CP-element group 346: 	 branch_block_stmt_655/lorx_xlhsx_xfalse697_ifx_xthen707_PhiReq/$exit
      -- 
    else_choice_transition_6015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2440_branch_ack_0, ack => zeropad3D_CP_2067_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	990 
    -- CP-element group 347: successors 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_Sample/ra
      -- 
    ra_6029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_0, ack => zeropad3D_CP_2067_elements(347)); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	990 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_Update/ca
      -- 
    ca_6034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_1, ack => zeropad3D_CP_2067_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	990 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_Sample/ra
      -- 
    ra_6043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2455_inst_ack_0, ack => zeropad3D_CP_2067_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	990 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_Update/ca
      -- 
    ca_6048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2455_inst_ack_1, ack => zeropad3D_CP_2067_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_Sample/rr
      -- 
    rr_6056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(351), ack => type_cast_2489_inst_req_0); -- 
    zeropad3D_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(348) & zeropad3D_CP_2067_elements(350);
      gj_zeropad3D_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_Sample/ra
      -- 
    ra_6057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2489_inst_ack_0, ack => zeropad3D_CP_2067_elements(352)); -- 
    -- CP-element group 353:  transition  input  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	990 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (16) 
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_Update/ca
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_resized_1
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_scaled_1
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_computed_1
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_resize_1/$entry
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_resize_1/$exit
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_resize_1/index_resize_req
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_resize_1/index_resize_ack
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_scale_1/$entry
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_scale_1/$exit
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_scale_1/scale_rename_req
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_index_scale_1/scale_rename_ack
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_Sample/req
      -- 
    ca_6062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2489_inst_ack_1, ack => zeropad3D_CP_2067_elements(353)); -- 
    req_6087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(353), ack => array_obj_ref_2495_index_offset_req_0); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	360 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_sample_complete
      -- CP-element group 354: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_Sample/ack
      -- 
    ack_6088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2495_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(354)); -- 
    -- CP-element group 355:  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	990 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (11) 
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_root_address_calculated
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_offset_calculated
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_Update/ack
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_base_plus_offset/$entry
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_base_plus_offset/$exit
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_base_plus_offset/sum_rename_req
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_base_plus_offset/sum_rename_ack
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_request/$entry
      -- CP-element group 355: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_request/req
      -- 
    ack_6093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2495_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(355)); -- 
    req_6102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(355), ack => addr_of_2496_final_reg_req_0); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_request/$exit
      -- CP-element group 356: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_request/ack
      -- 
    ack_6103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2496_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(356)); -- 
    -- CP-element group 357:  join  fork  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	990 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (28) 
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_complete/$exit
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_complete/ack
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_word_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_root_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_address_resized
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_addr_resize/$entry
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_addr_resize/$exit
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_addr_resize/base_resize_req
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_addr_resize/base_resize_ack
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_plus_offset/$entry
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_plus_offset/$exit
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_plus_offset/sum_rename_req
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_base_plus_offset/sum_rename_ack
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_word_addrgen/$entry
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_word_addrgen/$exit
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_word_addrgen/root_register_req
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_word_addrgen/root_register_ack
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/ptr_deref_2499_Split/$entry
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/ptr_deref_2499_Split/$exit
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/ptr_deref_2499_Split/split_req
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/ptr_deref_2499_Split/split_ack
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/word_access_start/$entry
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/word_access_start/word_0/$entry
      -- CP-element group 357: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/word_access_start/word_0/rr
      -- 
    ack_6108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2496_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(357)); -- 
    rr_6146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(357), ack => ptr_deref_2499_store_0_req_0); -- 
    -- CP-element group 358:  transition  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358:  members (5) 
      -- CP-element group 358: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_sample_completed_
      -- CP-element group 358: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/word_access_start/$exit
      -- CP-element group 358: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/word_access_start/word_0/$exit
      -- CP-element group 358: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Sample/word_access_start/word_0/ra
      -- 
    ra_6147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_store_0_ack_0, ack => zeropad3D_CP_2067_elements(358)); -- 
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	990 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (5) 
      -- CP-element group 359: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_update_completed_
      -- CP-element group 359: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Update/word_access_complete/$exit
      -- CP-element group 359: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Update/word_access_complete/word_0/$exit
      -- CP-element group 359: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Update/word_access_complete/word_0/ca
      -- 
    ca_6158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_store_0_ack_1, ack => zeropad3D_CP_2067_elements(359)); -- 
    -- CP-element group 360:  join  transition  place  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	354 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	991 
    -- CP-element group 360:  members (5) 
      -- CP-element group 360: 	 branch_block_stmt_655/ifx_xthen707_ifx_xend776
      -- CP-element group 360: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502__exit__
      -- CP-element group 360: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/$exit
      -- CP-element group 360: 	 branch_block_stmt_655/ifx_xthen707_ifx_xend776_PhiReq/$entry
      -- CP-element group 360: 	 branch_block_stmt_655/ifx_xthen707_ifx_xend776_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_360: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_360"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(354) & zeropad3D_CP_2067_elements(359);
      gj_zeropad3D_cp_element_group_360 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(360), clk => clk, reset => reset); --
    end block;
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	345 
    -- CP-element group 361: successors 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_Sample/ra
      -- 
    ra_6170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_0, ack => zeropad3D_CP_2067_elements(361)); -- 
    -- CP-element group 362:  fork  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	345 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362: 	371 
    -- CP-element group 362:  members (9) 
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2508_Update/ca
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_Sample/rr
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_Sample/rr
      -- 
    ca_6175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_1, ack => zeropad3D_CP_2067_elements(362)); -- 
    rr_6183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(362), ack => type_cast_2572_inst_req_0); -- 
    rr_6293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(362), ack => type_cast_2597_inst_req_0); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_Sample/ra
      -- 
    ra_6184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2572_inst_ack_0, ack => zeropad3D_CP_2067_elements(363)); -- 
    -- CP-element group 364:  transition  input  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	345 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (16) 
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2572_Update/ca
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_resized_1
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_scaled_1
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_computed_1
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_resize_1/$entry
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_resize_1/$exit
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_resize_1/index_resize_req
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_resize_1/index_resize_ack
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_scale_1/$entry
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_scale_1/$exit
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_scale_1/scale_rename_req
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_index_scale_1/scale_rename_ack
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_Sample/$entry
      -- CP-element group 364: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_Sample/req
      -- 
    ca_6189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2572_inst_ack_1, ack => zeropad3D_CP_2067_elements(364)); -- 
    req_6214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(364), ack => array_obj_ref_2578_index_offset_req_0); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	380 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_sample_complete
      -- CP-element group 365: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_Sample/ack
      -- 
    ack_6215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2578_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(365)); -- 
    -- CP-element group 366:  transition  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	345 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (11) 
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_root_address_calculated
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_offset_calculated
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_final_index_sum_regn_Update/ack
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_base_plus_offset/$entry
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_base_plus_offset/$exit
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_base_plus_offset/sum_rename_req
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2578_base_plus_offset/sum_rename_ack
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_request/$entry
      -- CP-element group 366: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_request/req
      -- 
    ack_6220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2578_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(366)); -- 
    req_6229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(366), ack => addr_of_2579_final_reg_req_0); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_request/$exit
      -- CP-element group 367: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_request/ack
      -- 
    ack_6230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2579_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(367)); -- 
    -- CP-element group 368:  join  fork  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	345 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (24) 
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_complete/$exit
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2579_complete/ack
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_sample_start_
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_address_calculated
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_word_address_calculated
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_root_address_calculated
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_address_resized
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_addr_resize/$entry
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_addr_resize/$exit
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_addr_resize/base_resize_req
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_addr_resize/base_resize_ack
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_plus_offset/$entry
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_plus_offset/$exit
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_plus_offset/sum_rename_req
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_base_plus_offset/sum_rename_ack
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_word_addrgen/$entry
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_word_addrgen/$exit
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_word_addrgen/root_register_req
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_word_addrgen/root_register_ack
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Sample/word_access_start/$entry
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Sample/word_access_start/word_0/$entry
      -- CP-element group 368: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Sample/word_access_start/word_0/rr
      -- 
    ack_6235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2579_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(368)); -- 
    rr_6268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(368), ack => ptr_deref_2583_load_0_req_0); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369:  members (5) 
      -- CP-element group 369: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Sample/word_access_start/$exit
      -- CP-element group 369: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Sample/word_access_start/word_0/$exit
      -- CP-element group 369: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Sample/word_access_start/word_0/ra
      -- 
    ra_6269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2583_load_0_ack_0, ack => zeropad3D_CP_2067_elements(369)); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	345 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	377 
    -- CP-element group 370:  members (9) 
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/word_access_complete/$exit
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/word_access_complete/word_0/$exit
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/word_access_complete/word_0/ca
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/ptr_deref_2583_Merge/$entry
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/ptr_deref_2583_Merge/$exit
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/ptr_deref_2583_Merge/merge_req
      -- CP-element group 370: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2583_Update/ptr_deref_2583_Merge/merge_ack
      -- 
    ca_6280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2583_load_0_ack_1, ack => zeropad3D_CP_2067_elements(370)); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	362 
    -- CP-element group 371: successors 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_Sample/ra
      -- 
    ra_6294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2597_inst_ack_0, ack => zeropad3D_CP_2067_elements(371)); -- 
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	345 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (16) 
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/type_cast_2597_Update/ca
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_resized_1
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_scaled_1
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_computed_1
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_resize_1/$entry
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_resize_1/$exit
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_resize_1/index_resize_req
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_resize_1/index_resize_ack
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_scale_1/$entry
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_scale_1/$exit
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_scale_1/scale_rename_req
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_index_scale_1/scale_rename_ack
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_Sample/req
      -- 
    ca_6299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2597_inst_ack_1, ack => zeropad3D_CP_2067_elements(372)); -- 
    req_6324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(372), ack => array_obj_ref_2603_index_offset_req_0); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	380 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_sample_complete
      -- CP-element group 373: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_Sample/$exit
      -- CP-element group 373: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_Sample/ack
      -- 
    ack_6325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2603_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(373)); -- 
    -- CP-element group 374:  transition  input  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	345 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (11) 
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_root_address_calculated
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_offset_calculated
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_Update/$exit
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_final_index_sum_regn_Update/ack
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_base_plus_offset/$entry
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_base_plus_offset/$exit
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_base_plus_offset/sum_rename_req
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/array_obj_ref_2603_base_plus_offset/sum_rename_ack
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_request/$entry
      -- CP-element group 374: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_request/req
      -- 
    ack_6330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2603_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(374)); -- 
    req_6339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(374), ack => addr_of_2604_final_reg_req_0); -- 
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_request/$exit
      -- CP-element group 375: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_request/ack
      -- 
    ack_6340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2604_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(375)); -- 
    -- CP-element group 376:  fork  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	345 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (19) 
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_complete/$exit
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/addr_of_2604_complete/ack
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_word_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_root_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_address_resized
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_addr_resize/$entry
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_addr_resize/$exit
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_addr_resize/base_resize_req
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_addr_resize/base_resize_ack
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_plus_offset/$entry
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_plus_offset/$exit
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_plus_offset/sum_rename_req
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_base_plus_offset/sum_rename_ack
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_word_addrgen/$entry
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_word_addrgen/$exit
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_word_addrgen/root_register_req
      -- CP-element group 376: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_word_addrgen/root_register_ack
      -- 
    ack_6345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2604_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	370 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (9) 
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/ptr_deref_2607_Split/$entry
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/ptr_deref_2607_Split/$exit
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/ptr_deref_2607_Split/split_req
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/ptr_deref_2607_Split/split_ack
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/word_access_start/$entry
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/word_access_start/word_0/$entry
      -- CP-element group 377: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/word_access_start/word_0/rr
      -- 
    rr_6383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(377), ack => ptr_deref_2607_store_0_req_0); -- 
    zeropad3D_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(370) & zeropad3D_CP_2067_elements(376);
      gj_zeropad3D_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378:  members (5) 
      -- CP-element group 378: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/word_access_start/$exit
      -- CP-element group 378: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/word_access_start/word_0/$exit
      -- CP-element group 378: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Sample/word_access_start/word_0/ra
      -- 
    ra_6384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2607_store_0_ack_0, ack => zeropad3D_CP_2067_elements(378)); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	345 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (5) 
      -- CP-element group 379: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Update/word_access_complete/$exit
      -- CP-element group 379: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Update/word_access_complete/word_0/$exit
      -- CP-element group 379: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/ptr_deref_2607_Update/word_access_complete/word_0/ca
      -- 
    ca_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2607_store_0_ack_1, ack => zeropad3D_CP_2067_elements(379)); -- 
    -- CP-element group 380:  join  transition  place  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	365 
    -- CP-element group 380: 	373 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	991 
    -- CP-element group 380:  members (5) 
      -- CP-element group 380: 	 branch_block_stmt_655/ifx_xelse728_ifx_xend776
      -- CP-element group 380: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609__exit__
      -- CP-element group 380: 	 branch_block_stmt_655/assign_stmt_2509_to_assign_stmt_2609/$exit
      -- CP-element group 380: 	 branch_block_stmt_655/ifx_xelse728_ifx_xend776_PhiReq/$entry
      -- CP-element group 380: 	 branch_block_stmt_655/ifx_xelse728_ifx_xend776_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(365) & zeropad3D_CP_2067_elements(373) & zeropad3D_CP_2067_elements(379);
      gj_zeropad3D_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	991 
    -- CP-element group 381: successors 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_Sample/ra
      -- 
    ra_6407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2615_inst_ack_0, ack => zeropad3D_CP_2067_elements(381)); -- 
    -- CP-element group 382:  branch  transition  place  input  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	991 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382: 	384 
    -- CP-element group 382:  members (13) 
      -- CP-element group 382: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629__exit__
      -- CP-element group 382: 	 branch_block_stmt_655/if_stmt_2630__entry__
      -- CP-element group 382: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/$exit
      -- CP-element group 382: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_Update/ca
      -- CP-element group 382: 	 branch_block_stmt_655/if_stmt_2630_dead_link/$entry
      -- CP-element group 382: 	 branch_block_stmt_655/if_stmt_2630_eval_test/$entry
      -- CP-element group 382: 	 branch_block_stmt_655/if_stmt_2630_eval_test/$exit
      -- CP-element group 382: 	 branch_block_stmt_655/if_stmt_2630_eval_test/branch_req
      -- CP-element group 382: 	 branch_block_stmt_655/R_cmp784_2631_place
      -- CP-element group 382: 	 branch_block_stmt_655/if_stmt_2630_if_link/$entry
      -- CP-element group 382: 	 branch_block_stmt_655/if_stmt_2630_else_link/$entry
      -- 
    ca_6412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2615_inst_ack_1, ack => zeropad3D_CP_2067_elements(382)); -- 
    branch_req_6420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(382), ack => if_stmt_2630_branch_req_0); -- 
    -- CP-element group 383:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	1000 
    -- CP-element group 383: 	1001 
    -- CP-element group 383: 	1003 
    -- CP-element group 383: 	1004 
    -- CP-element group 383: 	1006 
    -- CP-element group 383: 	1007 
    -- CP-element group 383:  members (40) 
      -- CP-element group 383: 	 branch_block_stmt_655/merge_stmt_2636__exit__
      -- CP-element group 383: 	 branch_block_stmt_655/assign_stmt_2642__entry__
      -- CP-element group 383: 	 branch_block_stmt_655/assign_stmt_2642__exit__
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827
      -- CP-element group 383: 	 branch_block_stmt_655/merge_stmt_2636_PhiReqMerge
      -- CP-element group 383: 	 branch_block_stmt_655/merge_stmt_2636_PhiAck/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/merge_stmt_2636_PhiAck/$exit
      -- CP-element group 383: 	 branch_block_stmt_655/merge_stmt_2636_PhiAck/dummy
      -- CP-element group 383: 	 branch_block_stmt_655/if_stmt_2630_if_link/$exit
      -- CP-element group 383: 	 branch_block_stmt_655/if_stmt_2630_if_link/if_choice_transition
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xend776_ifx_xthen786
      -- CP-element group 383: 	 branch_block_stmt_655/assign_stmt_2642/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/assign_stmt_2642/$exit
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xend776_ifx_xthen786_PhiReq/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xend776_ifx_xthen786_PhiReq/$exit
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Sample/rr
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Update/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Update/cr
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/Sample/rr
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/Update/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/Update/cr
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/Sample/rr
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/Update/$entry
      -- CP-element group 383: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2630_branch_ack_1, ack => zeropad3D_CP_2067_elements(383)); -- 
    rr_12210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(383), ack => type_cast_2726_inst_req_0); -- 
    cr_12215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(383), ack => type_cast_2726_inst_req_1); -- 
    rr_12233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(383), ack => type_cast_2733_inst_req_0); -- 
    cr_12238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(383), ack => type_cast_2733_inst_req_1); -- 
    rr_12256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(383), ack => type_cast_2739_inst_req_0); -- 
    cr_12261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(383), ack => type_cast_2739_inst_req_1); -- 
    -- CP-element group 384:  fork  transition  place  input  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	382 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384: 	386 
    -- CP-element group 384: 	387 
    -- CP-element group 384: 	388 
    -- CP-element group 384: 	390 
    -- CP-element group 384: 	393 
    -- CP-element group 384: 	395 
    -- CP-element group 384: 	396 
    -- CP-element group 384: 	397 
    -- CP-element group 384: 	399 
    -- CP-element group 384:  members (54) 
      -- CP-element group 384: 	 branch_block_stmt_655/merge_stmt_2644__exit__
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715__entry__
      -- CP-element group 384: 	 branch_block_stmt_655/if_stmt_2630_else_link/$exit
      -- CP-element group 384: 	 branch_block_stmt_655/if_stmt_2630_else_link/else_choice_transition
      -- CP-element group 384: 	 branch_block_stmt_655/ifx_xend776_ifx_xelse791
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_update_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_Sample/rr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_update_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_word_address_calculated
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_root_address_calculated
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Sample/word_access_start/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Sample/word_access_start/word_0/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Sample/word_access_start/word_0/rr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/word_access_complete/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/word_access_complete/word_0/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/word_access_complete/word_0/cr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_update_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_update_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_update_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_update_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_word_address_calculated
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_root_address_calculated
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Sample/word_access_start/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Sample/word_access_start/word_0/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Sample/word_access_start/word_0/rr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/word_access_complete/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/word_access_complete/word_0/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/word_access_complete/word_0/cr
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_update_start_
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_655/ifx_xend776_ifx_xelse791_PhiReq/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/ifx_xend776_ifx_xelse791_PhiReq/$exit
      -- CP-element group 384: 	 branch_block_stmt_655/merge_stmt_2644_PhiReqMerge
      -- CP-element group 384: 	 branch_block_stmt_655/merge_stmt_2644_PhiAck/$entry
      -- CP-element group 384: 	 branch_block_stmt_655/merge_stmt_2644_PhiAck/$exit
      -- CP-element group 384: 	 branch_block_stmt_655/merge_stmt_2644_PhiAck/dummy
      -- 
    else_choice_transition_6429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2630_branch_ack_0, ack => zeropad3D_CP_2067_elements(384)); -- 
    rr_6445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => type_cast_2654_inst_req_0); -- 
    cr_6450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => type_cast_2654_inst_req_1); -- 
    rr_6467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => LOAD_col_high_2657_load_0_req_0); -- 
    cr_6478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => LOAD_col_high_2657_load_0_req_1); -- 
    cr_6497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => type_cast_2661_inst_req_1); -- 
    cr_6511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => type_cast_2675_inst_req_1); -- 
    cr_6525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => type_cast_2691_inst_req_1); -- 
    rr_6542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => LOAD_row_high_2694_load_0_req_0); -- 
    cr_6553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => LOAD_row_high_2694_load_0_req_1); -- 
    cr_6572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(384), ack => type_cast_2698_inst_req_1); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_sample_completed_
      -- CP-element group 385: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_Sample/ra
      -- 
    ra_6446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2654_inst_ack_0, ack => zeropad3D_CP_2067_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	391 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_update_completed_
      -- CP-element group 386: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2654_Update/ca
      -- 
    ca_6451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2654_inst_ack_1, ack => zeropad3D_CP_2067_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	384 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (5) 
      -- CP-element group 387: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_sample_completed_
      -- CP-element group 387: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Sample/word_access_start/$exit
      -- CP-element group 387: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Sample/word_access_start/word_0/$exit
      -- CP-element group 387: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Sample/word_access_start/word_0/ra
      -- 
    ra_6468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2657_load_0_ack_0, ack => zeropad3D_CP_2067_elements(387)); -- 
    -- CP-element group 388:  transition  input  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	384 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (12) 
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/$exit
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/word_access_complete/$exit
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/word_access_complete/word_0/$exit
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/word_access_complete/word_0/ca
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/LOAD_col_high_2657_Merge/$entry
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/LOAD_col_high_2657_Merge/$exit
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/LOAD_col_high_2657_Merge/merge_req
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_col_high_2657_Update/LOAD_col_high_2657_Merge/merge_ack
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_sample_start_
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_Sample/$entry
      -- CP-element group 388: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_Sample/rr
      -- 
    ca_6479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2657_load_0_ack_1, ack => zeropad3D_CP_2067_elements(388)); -- 
    rr_6492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(388), ack => type_cast_2661_inst_req_0); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_sample_completed_
      -- CP-element group 389: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_Sample/ra
      -- 
    ra_6493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2661_inst_ack_0, ack => zeropad3D_CP_2067_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	384 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_update_completed_
      -- CP-element group 390: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2661_Update/ca
      -- 
    ca_6498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2661_inst_ack_1, ack => zeropad3D_CP_2067_elements(390)); -- 
    -- CP-element group 391:  join  transition  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	386 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_Sample/$entry
      -- CP-element group 391: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_Sample/rr
      -- 
    rr_6506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(391), ack => type_cast_2675_inst_req_0); -- 
    zeropad3D_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(386) & zeropad3D_CP_2067_elements(390);
      gj_zeropad3D_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_Sample/ra
      -- 
    ra_6507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2675_inst_ack_0, ack => zeropad3D_CP_2067_elements(392)); -- 
    -- CP-element group 393:  transition  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	384 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (6) 
      -- CP-element group 393: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2675_Update/ca
      -- CP-element group 393: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_Sample/rr
      -- 
    ca_6512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2675_inst_ack_1, ack => zeropad3D_CP_2067_elements(393)); -- 
    rr_6520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(393), ack => type_cast_2691_inst_req_0); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_Sample/ra
      -- 
    ra_6521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2691_inst_ack_0, ack => zeropad3D_CP_2067_elements(394)); -- 
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	384 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	400 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_update_completed_
      -- CP-element group 395: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2691_Update/ca
      -- 
    ca_6526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2691_inst_ack_1, ack => zeropad3D_CP_2067_elements(395)); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	384 
    -- CP-element group 396: successors 
    -- CP-element group 396:  members (5) 
      -- CP-element group 396: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_sample_completed_
      -- CP-element group 396: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Sample/word_access_start/$exit
      -- CP-element group 396: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Sample/word_access_start/word_0/$exit
      -- CP-element group 396: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Sample/word_access_start/word_0/ra
      -- 
    ra_6543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2694_load_0_ack_0, ack => zeropad3D_CP_2067_elements(396)); -- 
    -- CP-element group 397:  transition  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	384 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (12) 
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_update_completed_
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/word_access_complete/$exit
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/word_access_complete/word_0/$exit
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/word_access_complete/word_0/ca
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/LOAD_row_high_2694_Merge/$entry
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/LOAD_row_high_2694_Merge/$exit
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/LOAD_row_high_2694_Merge/merge_req
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/LOAD_row_high_2694_Update/LOAD_row_high_2694_Merge/merge_ack
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_Sample/rr
      -- 
    ca_6554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2694_load_0_ack_1, ack => zeropad3D_CP_2067_elements(397)); -- 
    rr_6567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(397), ack => type_cast_2698_inst_req_0); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_Sample/$exit
      -- CP-element group 398: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_Sample/ra
      -- 
    ra_6568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2698_inst_ack_0, ack => zeropad3D_CP_2067_elements(398)); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	384 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_Update/$exit
      -- CP-element group 399: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/type_cast_2698_Update/ca
      -- 
    ca_6573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2698_inst_ack_1, ack => zeropad3D_CP_2067_elements(399)); -- 
    -- CP-element group 400:  branch  join  transition  place  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	395 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400: 	402 
    -- CP-element group 400:  members (10) 
      -- CP-element group 400: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715__exit__
      -- CP-element group 400: 	 branch_block_stmt_655/if_stmt_2716__entry__
      -- CP-element group 400: 	 branch_block_stmt_655/assign_stmt_2650_to_assign_stmt_2715/$exit
      -- CP-element group 400: 	 branch_block_stmt_655/if_stmt_2716_dead_link/$entry
      -- CP-element group 400: 	 branch_block_stmt_655/if_stmt_2716_eval_test/$entry
      -- CP-element group 400: 	 branch_block_stmt_655/if_stmt_2716_eval_test/$exit
      -- CP-element group 400: 	 branch_block_stmt_655/if_stmt_2716_eval_test/branch_req
      -- CP-element group 400: 	 branch_block_stmt_655/R_cmp818_2717_place
      -- CP-element group 400: 	 branch_block_stmt_655/if_stmt_2716_if_link/$entry
      -- CP-element group 400: 	 branch_block_stmt_655/if_stmt_2716_else_link/$entry
      -- 
    branch_req_6581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(400), ack => if_stmt_2716_branch_req_0); -- 
    zeropad3D_cp_element_group_400: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_400"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(395) & zeropad3D_CP_2067_elements(399);
      gj_zeropad3D_cp_element_group_400 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(400), clk => clk, reset => reset); --
    end block;
    -- CP-element group 401:  fork  transition  place  input  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	1015 
    -- CP-element group 401: 	1016 
    -- CP-element group 401: 	1018 
    -- CP-element group 401: 	1019 
    -- CP-element group 401:  members (20) 
      -- CP-element group 401: 	 branch_block_stmt_655/if_stmt_2716_if_link/$exit
      -- CP-element group 401: 	 branch_block_stmt_655/if_stmt_2716_if_link/if_choice_transition
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/Sample/rr
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/Update/cr
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/Sample/rr
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2716_branch_ack_1, ack => zeropad3D_CP_2067_elements(401)); -- 
    rr_12289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(401), ack => type_cast_2748_inst_req_0); -- 
    cr_12294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(401), ack => type_cast_2748_inst_req_1); -- 
    rr_12312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(401), ack => type_cast_2752_inst_req_0); -- 
    cr_12317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(401), ack => type_cast_2752_inst_req_1); -- 
    -- CP-element group 402:  fork  transition  place  input  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	400 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	992 
    -- CP-element group 402: 	993 
    -- CP-element group 402: 	994 
    -- CP-element group 402: 	996 
    -- CP-element group 402: 	997 
    -- CP-element group 402:  members (22) 
      -- CP-element group 402: 	 branch_block_stmt_655/if_stmt_2716_else_link/$exit
      -- CP-element group 402: 	 branch_block_stmt_655/if_stmt_2716_else_link/else_choice_transition
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2723/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/Sample/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/Sample/rr
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/Update/cr
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/Sample/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/Sample/rr
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2716_branch_ack_0, ack => zeropad3D_CP_2067_elements(402)); -- 
    rr_12161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(402), ack => type_cast_2735_inst_req_0); -- 
    cr_12166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(402), ack => type_cast_2735_inst_req_1); -- 
    rr_12184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(402), ack => type_cast_2741_inst_req_0); -- 
    cr_12189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(402), ack => type_cast_2741_inst_req_1); -- 
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	1024 
    -- CP-element group 403: successors 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_sample_completed_
      -- CP-element group 403: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_Sample/ra
      -- 
    ra_6604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2756_inst_ack_0, ack => zeropad3D_CP_2067_elements(403)); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	1024 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	423 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_update_completed_
      -- CP-element group 404: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_Update/ca
      -- 
    ca_6609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2756_inst_ack_1, ack => zeropad3D_CP_2067_elements(404)); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	1024 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (5) 
      -- CP-element group 405: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_sample_completed_
      -- CP-element group 405: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Sample/$exit
      -- CP-element group 405: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Sample/word_access_start/$exit
      -- CP-element group 405: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Sample/word_access_start/word_0/$exit
      -- CP-element group 405: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Sample/word_access_start/word_0/ra
      -- 
    ra_6626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2765_load_0_ack_0, ack => zeropad3D_CP_2067_elements(405)); -- 
    -- CP-element group 406:  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	1024 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	419 
    -- CP-element group 406:  members (12) 
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/word_access_complete/word_0/ca
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/LOAD_pad_2765_Merge/$entry
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/LOAD_pad_2765_Merge/$exit
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/LOAD_pad_2765_Merge/merge_req
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/LOAD_pad_2765_Merge/merge_ack
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/word_access_complete/word_0/$exit
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/word_access_complete/$exit
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/$exit
      -- CP-element group 406: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_update_completed_
      -- 
    ca_6637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2765_load_0_ack_1, ack => zeropad3D_CP_2067_elements(406)); -- 
    rr_6791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(406), ack => type_cast_2795_inst_req_0); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	1024 
    -- CP-element group 407: successors 
    -- CP-element group 407:  members (5) 
      -- CP-element group 407: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_sample_completed_
      -- CP-element group 407: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Sample/word_access_start/word_0/ra
      -- CP-element group 407: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Sample/word_access_start/word_0/$exit
      -- CP-element group 407: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Sample/word_access_start/$exit
      -- 
    ra_6659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_2768_load_0_ack_0, ack => zeropad3D_CP_2067_elements(407)); -- 
    -- CP-element group 408:  transition  input  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	1024 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	413 
    -- CP-element group 408:  members (12) 
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_update_completed_
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/LOAD_depth_high_2768_Merge/merge_ack
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/LOAD_depth_high_2768_Merge/merge_req
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/LOAD_depth_high_2768_Merge/$exit
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/LOAD_depth_high_2768_Merge/$entry
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/word_access_complete/word_0/ca
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/word_access_complete/word_0/$exit
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/word_access_complete/$exit
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_Sample/rr
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_sample_start_
      -- 
    ca_6670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_2768_load_0_ack_1, ack => zeropad3D_CP_2067_elements(408)); -- 
    rr_6749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(408), ack => type_cast_2778_inst_req_0); -- 
    -- CP-element group 409:  transition  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	1024 
    -- CP-element group 409: successors 
    -- CP-element group 409:  members (5) 
      -- CP-element group 409: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Sample/word_access_start/$exit
      -- CP-element group 409: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Sample/word_access_start/word_0/$exit
      -- CP-element group 409: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Sample/word_access_start/word_0/ra
      -- CP-element group 409: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_sample_completed_
      -- 
    ra_6692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_2771_load_0_ack_0, ack => zeropad3D_CP_2067_elements(409)); -- 
    -- CP-element group 410:  fork  transition  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	1024 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	415 
    -- CP-element group 410: 	421 
    -- CP-element group 410:  members (15) 
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/word_access_complete/word_0/$exit
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/word_access_complete/word_0/ca
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/LOAD_out_depth_high_2771_Merge/$entry
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/LOAD_out_depth_high_2771_Merge/$exit
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/LOAD_out_depth_high_2771_Merge/merge_req
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/LOAD_out_depth_high_2771_Merge/merge_ack
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_sample_start_
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_Sample/$entry
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_Sample/rr
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/word_access_complete/$exit
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_update_completed_
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_Sample/rr
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_Sample/$entry
      -- CP-element group 410: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_sample_start_
      -- 
    ca_6703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_2771_load_0_ack_1, ack => zeropad3D_CP_2067_elements(410)); -- 
    rr_6763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(410), ack => type_cast_2782_inst_req_0); -- 
    rr_6805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(410), ack => type_cast_2799_inst_req_0); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	1024 
    -- CP-element group 411: successors 
    -- CP-element group 411:  members (5) 
      -- CP-element group 411: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_sample_completed_
      -- CP-element group 411: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Sample/$exit
      -- CP-element group 411: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Sample/word_access_start/word_0/ra
      -- CP-element group 411: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Sample/word_access_start/word_0/$exit
      -- CP-element group 411: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Sample/word_access_start/$exit
      -- 
    ra_6725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_2774_load_0_ack_0, ack => zeropad3D_CP_2067_elements(411)); -- 
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	1024 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	417 
    -- CP-element group 412:  members (12) 
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/$exit
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/word_access_complete/$exit
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/word_access_complete/word_0/$exit
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_update_completed_
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/word_access_complete/word_0/ca
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/LOAD_out_col_high_2774_Merge/$entry
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_Sample/rr
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_Sample/$entry
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_sample_start_
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/LOAD_out_col_high_2774_Merge/merge_ack
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/LOAD_out_col_high_2774_Merge/merge_req
      -- CP-element group 412: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/LOAD_out_col_high_2774_Merge/$exit
      -- 
    ca_6736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_2774_load_0_ack_1, ack => zeropad3D_CP_2067_elements(412)); -- 
    rr_6777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(412), ack => type_cast_2786_inst_req_0); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	408 
    -- CP-element group 413: successors 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_Sample/ra
      -- CP-element group 413: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_Sample/$exit
      -- CP-element group 413: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_sample_completed_
      -- 
    ra_6750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2778_inst_ack_0, ack => zeropad3D_CP_2067_elements(413)); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	1024 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	423 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_Update/ca
      -- CP-element group 414: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_Update/$exit
      -- CP-element group 414: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_update_completed_
      -- 
    ca_6755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2778_inst_ack_1, ack => zeropad3D_CP_2067_elements(414)); -- 
    -- CP-element group 415:  transition  input  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	410 
    -- CP-element group 415: successors 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_Sample/ra
      -- CP-element group 415: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_sample_completed_
      -- 
    ra_6764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2782_inst_ack_0, ack => zeropad3D_CP_2067_elements(415)); -- 
    -- CP-element group 416:  transition  input  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	1024 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	423 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_Update/ca
      -- CP-element group 416: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_update_completed_
      -- 
    ca_6769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2782_inst_ack_1, ack => zeropad3D_CP_2067_elements(416)); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	412 
    -- CP-element group 417: successors 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_Sample/ra
      -- CP-element group 417: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_Sample/$exit
      -- CP-element group 417: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_sample_completed_
      -- 
    ra_6778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2786_inst_ack_0, ack => zeropad3D_CP_2067_elements(417)); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	1024 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	423 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_Update/ca
      -- CP-element group 418: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_Update/$exit
      -- CP-element group 418: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_update_completed_
      -- 
    ca_6783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2786_inst_ack_1, ack => zeropad3D_CP_2067_elements(418)); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	406 
    -- CP-element group 419: successors 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_sample_completed_
      -- CP-element group 419: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_Sample/ra
      -- 
    ra_6792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2795_inst_ack_0, ack => zeropad3D_CP_2067_elements(419)); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	1024 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	423 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_Update/ca
      -- 
    ca_6797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2795_inst_ack_1, ack => zeropad3D_CP_2067_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	410 
    -- CP-element group 421: successors 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_sample_completed_
      -- CP-element group 421: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_Sample/$exit
      -- CP-element group 421: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_Sample/ra
      -- 
    ra_6806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2799_inst_ack_0, ack => zeropad3D_CP_2067_elements(421)); -- 
    -- CP-element group 422:  transition  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	1024 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_update_completed_
      -- CP-element group 422: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_Update/$exit
      -- CP-element group 422: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_Update/ca
      -- 
    ca_6811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2799_inst_ack_1, ack => zeropad3D_CP_2067_elements(422)); -- 
    -- CP-element group 423:  join  fork  transition  place  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	404 
    -- CP-element group 423: 	414 
    -- CP-element group 423: 	416 
    -- CP-element group 423: 	418 
    -- CP-element group 423: 	420 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	1035 
    -- CP-element group 423: 	1036 
    -- CP-element group 423: 	1037 
    -- CP-element group 423: 	1039 
    -- CP-element group 423:  members (16) 
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888
      -- CP-element group 423: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841__exit__
      -- CP-element group 423: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/$exit
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2844/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/Sample/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/Sample/rr
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/Update/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/Update/cr
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2857/$entry
      -- CP-element group 423: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/$entry
      -- 
    rr_12424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(423), ack => type_cast_2854_inst_req_0); -- 
    cr_12429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(423), ack => type_cast_2854_inst_req_1); -- 
    zeropad3D_cp_element_group_423: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_423"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(404) & zeropad3D_CP_2067_elements(414) & zeropad3D_CP_2067_elements(416) & zeropad3D_CP_2067_elements(418) & zeropad3D_CP_2067_elements(420) & zeropad3D_CP_2067_elements(422);
      gj_zeropad3D_cp_element_group_423 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 424:  transition  input  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	1045 
    -- CP-element group 424: successors 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_Sample/ra
      -- CP-element group 424: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_Sample/$exit
      -- CP-element group 424: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_sample_completed_
      -- 
    ra_6823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2868_inst_ack_0, ack => zeropad3D_CP_2067_elements(424)); -- 
    -- CP-element group 425:  branch  transition  place  input  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	1045 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425: 	427 
    -- CP-element group 425:  members (13) 
      -- CP-element group 425: 	 branch_block_stmt_655/if_stmt_2877__entry__
      -- CP-element group 425: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876__exit__
      -- CP-element group 425: 	 branch_block_stmt_655/if_stmt_2877_eval_test/$entry
      -- CP-element group 425: 	 branch_block_stmt_655/if_stmt_2877_eval_test/$exit
      -- CP-element group 425: 	 branch_block_stmt_655/if_stmt_2877_eval_test/branch_req
      -- CP-element group 425: 	 branch_block_stmt_655/if_stmt_2877_if_link/$entry
      -- CP-element group 425: 	 branch_block_stmt_655/if_stmt_2877_dead_link/$entry
      -- CP-element group 425: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_Update/ca
      -- CP-element group 425: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_Update/$exit
      -- CP-element group 425: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_update_completed_
      -- CP-element group 425: 	 branch_block_stmt_655/R_cmp893_2878_place
      -- CP-element group 425: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/$exit
      -- CP-element group 425: 	 branch_block_stmt_655/if_stmt_2877_else_link/$entry
      -- 
    ca_6828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2868_inst_ack_1, ack => zeropad3D_CP_2067_elements(425)); -- 
    branch_req_6836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(425), ack => if_stmt_2877_branch_req_0); -- 
    -- CP-element group 426:  transition  place  input  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	1046 
    -- CP-element group 426:  members (5) 
      -- CP-element group 426: 	 branch_block_stmt_655/whilex_xbody888_ifx_xthen925
      -- CP-element group 426: 	 branch_block_stmt_655/if_stmt_2877_if_link/if_choice_transition
      -- CP-element group 426: 	 branch_block_stmt_655/if_stmt_2877_if_link/$exit
      -- CP-element group 426: 	 branch_block_stmt_655/whilex_xbody888_ifx_xthen925_PhiReq/$entry
      -- CP-element group 426: 	 branch_block_stmt_655/whilex_xbody888_ifx_xthen925_PhiReq/$exit
      -- 
    if_choice_transition_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2877_branch_ack_1, ack => zeropad3D_CP_2067_elements(426)); -- 
    -- CP-element group 427:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	425 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427: 	429 
    -- CP-element group 427: 	431 
    -- CP-element group 427:  members (27) 
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914__entry__
      -- CP-element group 427: 	 branch_block_stmt_655/merge_stmt_2883__exit__
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_Update/cr
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_update_start_
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/word_access_complete/word_0/cr
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/word_access_complete/word_0/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/word_access_complete/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Sample/word_access_start/word_0/rr
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Sample/word_access_start/word_0/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Sample/word_access_start/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/whilex_xbody888_lorx_xlhsx_xfalse895
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_root_address_calculated
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_word_address_calculated
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_update_start_
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/if_stmt_2877_else_link/else_choice_transition
      -- CP-element group 427: 	 branch_block_stmt_655/if_stmt_2877_else_link/$exit
      -- CP-element group 427: 	 branch_block_stmt_655/whilex_xbody888_lorx_xlhsx_xfalse895_PhiReq/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/whilex_xbody888_lorx_xlhsx_xfalse895_PhiReq/$exit
      -- CP-element group 427: 	 branch_block_stmt_655/merge_stmt_2883_PhiReqMerge
      -- CP-element group 427: 	 branch_block_stmt_655/merge_stmt_2883_PhiAck/$entry
      -- CP-element group 427: 	 branch_block_stmt_655/merge_stmt_2883_PhiAck/$exit
      -- CP-element group 427: 	 branch_block_stmt_655/merge_stmt_2883_PhiAck/dummy
      -- 
    else_choice_transition_6845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2877_branch_ack_0, ack => zeropad3D_CP_2067_elements(427)); -- 
    cr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(427), ack => type_cast_2889_inst_req_1); -- 
    cr_6877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(427), ack => LOAD_row_high_2885_load_0_req_1); -- 
    rr_6866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(427), ack => LOAD_row_high_2885_load_0_req_0); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428:  members (5) 
      -- CP-element group 428: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Sample/word_access_start/word_0/ra
      -- CP-element group 428: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Sample/word_access_start/word_0/$exit
      -- CP-element group 428: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Sample/word_access_start/$exit
      -- CP-element group 428: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_sample_completed_
      -- 
    ra_6867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2885_load_0_ack_0, ack => zeropad3D_CP_2067_elements(428)); -- 
    -- CP-element group 429:  transition  input  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	427 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (12) 
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_sample_start_
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/LOAD_row_high_2885_Merge/merge_ack
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/LOAD_row_high_2885_Merge/merge_req
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/LOAD_row_high_2885_Merge/$exit
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/LOAD_row_high_2885_Merge/$entry
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/word_access_complete/word_0/ca
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/word_access_complete/word_0/$exit
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/word_access_complete/$exit
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/LOAD_row_high_2885_update_completed_
      -- 
    ca_6878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2885_load_0_ack_1, ack => zeropad3D_CP_2067_elements(429)); -- 
    rr_6891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(429), ack => type_cast_2889_inst_req_0); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_Sample/$exit
      -- CP-element group 430: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_Sample/ra
      -- CP-element group 430: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_sample_completed_
      -- 
    ra_6892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2889_inst_ack_0, ack => zeropad3D_CP_2067_elements(430)); -- 
    -- CP-element group 431:  branch  transition  place  input  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	427 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	432 
    -- CP-element group 431: 	433 
    -- CP-element group 431:  members (13) 
      -- CP-element group 431: 	 branch_block_stmt_655/if_stmt_2915__entry__
      -- CP-element group 431: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914__exit__
      -- CP-element group 431: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_update_completed_
      -- CP-element group 431: 	 branch_block_stmt_655/R_cmp905_2916_place
      -- CP-element group 431: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_Update/$exit
      -- CP-element group 431: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/type_cast_2889_Update/ca
      -- CP-element group 431: 	 branch_block_stmt_655/if_stmt_2915_else_link/$entry
      -- CP-element group 431: 	 branch_block_stmt_655/if_stmt_2915_if_link/$entry
      -- CP-element group 431: 	 branch_block_stmt_655/if_stmt_2915_eval_test/branch_req
      -- CP-element group 431: 	 branch_block_stmt_655/if_stmt_2915_eval_test/$exit
      -- CP-element group 431: 	 branch_block_stmt_655/if_stmt_2915_eval_test/$entry
      -- CP-element group 431: 	 branch_block_stmt_655/assign_stmt_2886_to_assign_stmt_2914/$exit
      -- CP-element group 431: 	 branch_block_stmt_655/if_stmt_2915_dead_link/$entry
      -- 
    ca_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2889_inst_ack_1, ack => zeropad3D_CP_2067_elements(431)); -- 
    branch_req_6905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(431), ack => if_stmt_2915_branch_req_0); -- 
    -- CP-element group 432:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	431 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	434 
    -- CP-element group 432: 	435 
    -- CP-element group 432:  members (18) 
      -- CP-element group 432: 	 branch_block_stmt_655/merge_stmt_2921__exit__
      -- CP-element group 432: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933__entry__
      -- CP-element group 432: 	 branch_block_stmt_655/lorx_xlhsx_xfalse895_lorx_xlhsx_xfalse907
      -- CP-element group 432: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_Update/cr
      -- CP-element group 432: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_Update/$entry
      -- CP-element group 432: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_Sample/rr
      -- CP-element group 432: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_Sample/$entry
      -- CP-element group 432: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_update_start_
      -- CP-element group 432: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_sample_start_
      -- CP-element group 432: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/$entry
      -- CP-element group 432: 	 branch_block_stmt_655/if_stmt_2915_if_link/if_choice_transition
      -- CP-element group 432: 	 branch_block_stmt_655/if_stmt_2915_if_link/$exit
      -- CP-element group 432: 	 branch_block_stmt_655/lorx_xlhsx_xfalse895_lorx_xlhsx_xfalse907_PhiReq/$entry
      -- CP-element group 432: 	 branch_block_stmt_655/lorx_xlhsx_xfalse895_lorx_xlhsx_xfalse907_PhiReq/$exit
      -- CP-element group 432: 	 branch_block_stmt_655/merge_stmt_2921_PhiReqMerge
      -- CP-element group 432: 	 branch_block_stmt_655/merge_stmt_2921_PhiAck/$entry
      -- CP-element group 432: 	 branch_block_stmt_655/merge_stmt_2921_PhiAck/$exit
      -- CP-element group 432: 	 branch_block_stmt_655/merge_stmt_2921_PhiAck/dummy
      -- 
    if_choice_transition_6910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2915_branch_ack_1, ack => zeropad3D_CP_2067_elements(432)); -- 
    cr_6932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(432), ack => type_cast_2925_inst_req_1); -- 
    rr_6927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(432), ack => type_cast_2925_inst_req_0); -- 
    -- CP-element group 433:  transition  place  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	431 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	1046 
    -- CP-element group 433:  members (5) 
      -- CP-element group 433: 	 branch_block_stmt_655/lorx_xlhsx_xfalse895_ifx_xthen925
      -- CP-element group 433: 	 branch_block_stmt_655/if_stmt_2915_else_link/else_choice_transition
      -- CP-element group 433: 	 branch_block_stmt_655/if_stmt_2915_else_link/$exit
      -- CP-element group 433: 	 branch_block_stmt_655/lorx_xlhsx_xfalse895_ifx_xthen925_PhiReq/$entry
      -- CP-element group 433: 	 branch_block_stmt_655/lorx_xlhsx_xfalse895_ifx_xthen925_PhiReq/$exit
      -- 
    else_choice_transition_6914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2915_branch_ack_0, ack => zeropad3D_CP_2067_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	432 
    -- CP-element group 434: successors 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_Sample/ra
      -- CP-element group 434: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_sample_completed_
      -- 
    ra_6928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2925_inst_ack_0, ack => zeropad3D_CP_2067_elements(434)); -- 
    -- CP-element group 435:  branch  transition  place  input  output  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	432 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435: 	437 
    -- CP-element group 435:  members (13) 
      -- CP-element group 435: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933__exit__
      -- CP-element group 435: 	 branch_block_stmt_655/if_stmt_2934__entry__
      -- CP-element group 435: 	 branch_block_stmt_655/R_cmp912_2935_place
      -- CP-element group 435: 	 branch_block_stmt_655/if_stmt_2934_else_link/$entry
      -- CP-element group 435: 	 branch_block_stmt_655/if_stmt_2934_if_link/$entry
      -- CP-element group 435: 	 branch_block_stmt_655/if_stmt_2934_eval_test/branch_req
      -- CP-element group 435: 	 branch_block_stmt_655/if_stmt_2934_eval_test/$exit
      -- CP-element group 435: 	 branch_block_stmt_655/if_stmt_2934_eval_test/$entry
      -- CP-element group 435: 	 branch_block_stmt_655/if_stmt_2934_dead_link/$entry
      -- CP-element group 435: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_Update/ca
      -- CP-element group 435: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/type_cast_2925_update_completed_
      -- CP-element group 435: 	 branch_block_stmt_655/assign_stmt_2926_to_assign_stmt_2933/$exit
      -- 
    ca_6933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2925_inst_ack_1, ack => zeropad3D_CP_2067_elements(435)); -- 
    branch_req_6941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(435), ack => if_stmt_2934_branch_req_0); -- 
    -- CP-element group 436:  transition  place  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	1046 
    -- CP-element group 436:  members (5) 
      -- CP-element group 436: 	 branch_block_stmt_655/lorx_xlhsx_xfalse907_ifx_xthen925
      -- CP-element group 436: 	 branch_block_stmt_655/if_stmt_2934_if_link/if_choice_transition
      -- CP-element group 436: 	 branch_block_stmt_655/if_stmt_2934_if_link/$exit
      -- CP-element group 436: 	 branch_block_stmt_655/lorx_xlhsx_xfalse907_ifx_xthen925_PhiReq/$entry
      -- CP-element group 436: 	 branch_block_stmt_655/lorx_xlhsx_xfalse907_ifx_xthen925_PhiReq/$exit
      -- 
    if_choice_transition_6946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2934_branch_ack_1, ack => zeropad3D_CP_2067_elements(436)); -- 
    -- CP-element group 437:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	435 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	438 
    -- CP-element group 437: 	439 
    -- CP-element group 437: 	441 
    -- CP-element group 437:  members (27) 
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965__entry__
      -- CP-element group 437: 	 branch_block_stmt_655/merge_stmt_2940__exit__
      -- CP-element group 437: 	 branch_block_stmt_655/if_stmt_2934_else_link/$exit
      -- CP-element group 437: 	 branch_block_stmt_655/if_stmt_2934_else_link/else_choice_transition
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_sample_start_
      -- CP-element group 437: 	 branch_block_stmt_655/lorx_xlhsx_xfalse907_lorx_xlhsx_xfalse914
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Sample/word_access_start/word_0/rr
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_update_start_
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Sample/word_access_start/word_0/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/word_access_complete/word_0/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_root_address_calculated
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/word_access_complete/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Sample/word_access_start/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_Update/cr
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_word_address_calculated
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_Update/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_update_start_
      -- CP-element group 437: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/word_access_complete/word_0/cr
      -- CP-element group 437: 	 branch_block_stmt_655/lorx_xlhsx_xfalse907_lorx_xlhsx_xfalse914_PhiReq/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/lorx_xlhsx_xfalse907_lorx_xlhsx_xfalse914_PhiReq/$exit
      -- CP-element group 437: 	 branch_block_stmt_655/merge_stmt_2940_PhiReqMerge
      -- CP-element group 437: 	 branch_block_stmt_655/merge_stmt_2940_PhiAck/$entry
      -- CP-element group 437: 	 branch_block_stmt_655/merge_stmt_2940_PhiAck/$exit
      -- CP-element group 437: 	 branch_block_stmt_655/merge_stmt_2940_PhiAck/dummy
      -- 
    else_choice_transition_6950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2934_branch_ack_0, ack => zeropad3D_CP_2067_elements(437)); -- 
    rr_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(437), ack => LOAD_col_high_2942_load_0_req_0); -- 
    cr_7001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(437), ack => type_cast_2946_inst_req_1); -- 
    cr_6982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(437), ack => LOAD_col_high_2942_load_0_req_1); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	437 
    -- CP-element group 438: successors 
    -- CP-element group 438:  members (5) 
      -- CP-element group 438: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Sample/word_access_start/word_0/$exit
      -- CP-element group 438: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_sample_completed_
      -- CP-element group 438: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Sample/word_access_start/word_0/ra
      -- CP-element group 438: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Sample/word_access_start/$exit
      -- 
    ra_6972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2942_load_0_ack_0, ack => zeropad3D_CP_2067_elements(438)); -- 
    -- CP-element group 439:  transition  input  output  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	437 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439:  members (12) 
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_update_completed_
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/LOAD_col_high_2942_Merge/$entry
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_Sample/rr
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_sample_start_
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/LOAD_col_high_2942_Merge/merge_ack
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/LOAD_col_high_2942_Merge/merge_req
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/LOAD_col_high_2942_Merge/$exit
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/word_access_complete/word_0/ca
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_Sample/$entry
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/word_access_complete/word_0/$exit
      -- CP-element group 439: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/LOAD_col_high_2942_Update/word_access_complete/$exit
      -- 
    ca_6983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2942_load_0_ack_1, ack => zeropad3D_CP_2067_elements(439)); -- 
    rr_6996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(439), ack => type_cast_2946_inst_req_0); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_Sample/ra
      -- CP-element group 440: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_Sample/$exit
      -- CP-element group 440: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_sample_completed_
      -- 
    ra_6997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2946_inst_ack_0, ack => zeropad3D_CP_2067_elements(440)); -- 
    -- CP-element group 441:  branch  transition  place  input  output  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	437 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441: 	443 
    -- CP-element group 441:  members (13) 
      -- CP-element group 441: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965__exit__
      -- CP-element group 441: 	 branch_block_stmt_655/if_stmt_2966__entry__
      -- CP-element group 441: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/$exit
      -- CP-element group 441: 	 branch_block_stmt_655/R_cmp923_2967_place
      -- CP-element group 441: 	 branch_block_stmt_655/if_stmt_2966_else_link/$entry
      -- CP-element group 441: 	 branch_block_stmt_655/if_stmt_2966_dead_link/$entry
      -- CP-element group 441: 	 branch_block_stmt_655/if_stmt_2966_if_link/$entry
      -- CP-element group 441: 	 branch_block_stmt_655/if_stmt_2966_eval_test/branch_req
      -- CP-element group 441: 	 branch_block_stmt_655/if_stmt_2966_eval_test/$exit
      -- CP-element group 441: 	 branch_block_stmt_655/if_stmt_2966_eval_test/$entry
      -- CP-element group 441: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_Update/ca
      -- CP-element group 441: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_Update/$exit
      -- CP-element group 441: 	 branch_block_stmt_655/assign_stmt_2943_to_assign_stmt_2965/type_cast_2946_update_completed_
      -- 
    ca_7002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2946_inst_ack_1, ack => zeropad3D_CP_2067_elements(441)); -- 
    branch_req_7010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(441), ack => if_stmt_2966_branch_req_0); -- 
    -- CP-element group 442:  fork  transition  place  input  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	441 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	458 
    -- CP-element group 442: 	459 
    -- CP-element group 442: 	461 
    -- CP-element group 442: 	463 
    -- CP-element group 442: 	465 
    -- CP-element group 442: 	467 
    -- CP-element group 442: 	469 
    -- CP-element group 442: 	471 
    -- CP-element group 442: 	473 
    -- CP-element group 442: 	476 
    -- CP-element group 442:  members (46) 
      -- CP-element group 442: 	 branch_block_stmt_655/merge_stmt_3030__exit__
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135__entry__
      -- CP-element group 442: 	 branch_block_stmt_655/lorx_xlhsx_xfalse914_ifx_xelse946
      -- CP-element group 442: 	 branch_block_stmt_655/if_stmt_2966_if_link/if_choice_transition
      -- CP-element group 442: 	 branch_block_stmt_655/if_stmt_2966_if_link/$exit
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_sample_start_
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_update_start_
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_Sample/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_Sample/rr
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_update_start_
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_update_start_
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_update_start
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_Update/req
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_complete/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_complete/req
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_update_start_
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/word_access_complete/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/word_access_complete/word_0/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/word_access_complete/word_0/cr
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_update_start_
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_Update/cr
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_update_start_
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_update_start
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_Update/req
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_complete/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_complete/req
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_update_start_
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Update/word_access_complete/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Update/word_access_complete/word_0/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Update/word_access_complete/word_0/cr
      -- CP-element group 442: 	 branch_block_stmt_655/lorx_xlhsx_xfalse914_ifx_xelse946_PhiReq/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/lorx_xlhsx_xfalse914_ifx_xelse946_PhiReq/$exit
      -- CP-element group 442: 	 branch_block_stmt_655/merge_stmt_3030_PhiReqMerge
      -- CP-element group 442: 	 branch_block_stmt_655/merge_stmt_3030_PhiAck/$entry
      -- CP-element group 442: 	 branch_block_stmt_655/merge_stmt_3030_PhiAck/$exit
      -- CP-element group 442: 	 branch_block_stmt_655/merge_stmt_3030_PhiAck/dummy
      -- 
    if_choice_transition_7015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2966_branch_ack_1, ack => zeropad3D_CP_2067_elements(442)); -- 
    rr_7173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => type_cast_3034_inst_req_0); -- 
    cr_7178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => type_cast_3034_inst_req_1); -- 
    cr_7192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => type_cast_3098_inst_req_1); -- 
    req_7223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => array_obj_ref_3104_index_offset_req_1); -- 
    req_7238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => addr_of_3105_final_reg_req_1); -- 
    cr_7283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => ptr_deref_3109_load_0_req_1); -- 
    cr_7302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => type_cast_3123_inst_req_1); -- 
    req_7333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => array_obj_ref_3129_index_offset_req_1); -- 
    req_7348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => addr_of_3130_final_reg_req_1); -- 
    cr_7398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(442), ack => ptr_deref_3133_store_0_req_1); -- 
    -- CP-element group 443:  transition  place  input  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	441 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	1046 
    -- CP-element group 443:  members (5) 
      -- CP-element group 443: 	 branch_block_stmt_655/if_stmt_2966_else_link/$exit
      -- CP-element group 443: 	 branch_block_stmt_655/if_stmt_2966_else_link/else_choice_transition
      -- CP-element group 443: 	 branch_block_stmt_655/lorx_xlhsx_xfalse914_ifx_xthen925
      -- CP-element group 443: 	 branch_block_stmt_655/lorx_xlhsx_xfalse914_ifx_xthen925_PhiReq/$entry
      -- CP-element group 443: 	 branch_block_stmt_655/lorx_xlhsx_xfalse914_ifx_xthen925_PhiReq/$exit
      -- 
    else_choice_transition_7019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2966_branch_ack_0, ack => zeropad3D_CP_2067_elements(443)); -- 
    -- CP-element group 444:  transition  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	1046 
    -- CP-element group 444: successors 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_sample_completed_
      -- CP-element group 444: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_Sample/ra
      -- CP-element group 444: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_Sample/$exit
      -- 
    ra_7033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2976_inst_ack_0, ack => zeropad3D_CP_2067_elements(444)); -- 
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	1046 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	448 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_Update/ca
      -- CP-element group 445: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_update_completed_
      -- 
    ca_7038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2976_inst_ack_1, ack => zeropad3D_CP_2067_elements(445)); -- 
    -- CP-element group 446:  transition  input  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	1046 
    -- CP-element group 446: successors 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_sample_completed_
      -- CP-element group 446: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_Sample/ra
      -- CP-element group 446: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_Sample/$exit
      -- 
    ra_7047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2981_inst_ack_0, ack => zeropad3D_CP_2067_elements(446)); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	1046 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_update_completed_
      -- CP-element group 447: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_Update/ca
      -- CP-element group 447: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_Update/$exit
      -- 
    ca_7052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2981_inst_ack_1, ack => zeropad3D_CP_2067_elements(447)); -- 
    -- CP-element group 448:  join  transition  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	445 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_Sample/rr
      -- CP-element group 448: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_Sample/$entry
      -- CP-element group 448: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_sample_start_
      -- 
    rr_7060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(448), ack => type_cast_3015_inst_req_0); -- 
    zeropad3D_cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(445) & zeropad3D_CP_2067_elements(447);
      gj_zeropad3D_cp_element_group_448 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 449:  transition  input  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_Sample/ra
      -- CP-element group 449: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_Sample/$exit
      -- CP-element group 449: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_sample_completed_
      -- 
    ra_7061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3015_inst_ack_0, ack => zeropad3D_CP_2067_elements(449)); -- 
    -- CP-element group 450:  transition  input  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	1046 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (16) 
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_Update/ca
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_Update/$exit
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_update_completed_
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_resized_1
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_scaled_1
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_computed_1
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_resize_1/$entry
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_resize_1/$exit
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_resize_1/index_resize_req
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_resize_1/index_resize_ack
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_scale_1/$entry
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_scale_1/$exit
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_scale_1/scale_rename_req
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_index_scale_1/scale_rename_ack
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_Sample/$entry
      -- CP-element group 450: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_Sample/req
      -- 
    ca_7066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3015_inst_ack_1, ack => zeropad3D_CP_2067_elements(450)); -- 
    req_7091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(450), ack => array_obj_ref_3021_index_offset_req_0); -- 
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	457 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_sample_complete
      -- CP-element group 451: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_Sample/$exit
      -- CP-element group 451: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_Sample/ack
      -- 
    ack_7092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3021_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(451)); -- 
    -- CP-element group 452:  transition  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	1046 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (11) 
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_root_address_calculated
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_offset_calculated
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_Update/$exit
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_Update/ack
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_base_plus_offset/$entry
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_base_plus_offset/$exit
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_base_plus_offset/sum_rename_req
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_base_plus_offset/sum_rename_ack
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_request/$entry
      -- CP-element group 452: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_request/req
      -- 
    ack_7097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3021_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(452)); -- 
    req_7106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(452), ack => addr_of_3022_final_reg_req_0); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_sample_completed_
      -- CP-element group 453: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_request/$exit
      -- CP-element group 453: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_request/ack
      -- 
    ack_7107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3022_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(453)); -- 
    -- CP-element group 454:  join  fork  transition  input  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	1046 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (28) 
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_update_completed_
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_complete/$exit
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_complete/ack
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_sample_start_
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_address_calculated
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_word_address_calculated
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_root_address_calculated
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_address_resized
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_addr_resize/$entry
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_addr_resize/$exit
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_addr_resize/base_resize_req
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_addr_resize/base_resize_ack
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_plus_offset/$entry
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_plus_offset/$exit
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_plus_offset/sum_rename_req
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_base_plus_offset/sum_rename_ack
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_word_addrgen/$entry
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_word_addrgen/$exit
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_word_addrgen/root_register_req
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_word_addrgen/root_register_ack
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/ptr_deref_3025_Split/$entry
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/ptr_deref_3025_Split/$exit
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/ptr_deref_3025_Split/split_req
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/ptr_deref_3025_Split/split_ack
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/word_access_start/$entry
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/word_access_start/word_0/$entry
      -- CP-element group 454: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/word_access_start/word_0/rr
      -- 
    ack_7112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3022_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(454)); -- 
    rr_7150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(454), ack => ptr_deref_3025_store_0_req_0); -- 
    -- CP-element group 455:  transition  input  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455:  members (5) 
      -- CP-element group 455: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_sample_completed_
      -- CP-element group 455: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/word_access_start/$exit
      -- CP-element group 455: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/word_access_start/word_0/$exit
      -- CP-element group 455: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Sample/word_access_start/word_0/ra
      -- 
    ra_7151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3025_store_0_ack_0, ack => zeropad3D_CP_2067_elements(455)); -- 
    -- CP-element group 456:  transition  input  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	1046 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (5) 
      -- CP-element group 456: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_update_completed_
      -- CP-element group 456: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Update/word_access_complete/$exit
      -- CP-element group 456: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Update/word_access_complete/word_0/$exit
      -- CP-element group 456: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Update/word_access_complete/word_0/ca
      -- 
    ca_7162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3025_store_0_ack_1, ack => zeropad3D_CP_2067_elements(456)); -- 
    -- CP-element group 457:  join  transition  place  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	451 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	1047 
    -- CP-element group 457:  members (5) 
      -- CP-element group 457: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028__exit__
      -- CP-element group 457: 	 branch_block_stmt_655/ifx_xthen925_ifx_xend994
      -- CP-element group 457: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/$exit
      -- CP-element group 457: 	 branch_block_stmt_655/ifx_xthen925_ifx_xend994_PhiReq/$entry
      -- CP-element group 457: 	 branch_block_stmt_655/ifx_xthen925_ifx_xend994_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(451) & zeropad3D_CP_2067_elements(456);
      gj_zeropad3D_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  transition  input  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	442 
    -- CP-element group 458: successors 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_sample_completed_
      -- CP-element group 458: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_Sample/$exit
      -- CP-element group 458: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_Sample/ra
      -- 
    ra_7174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3034_inst_ack_0, ack => zeropad3D_CP_2067_elements(458)); -- 
    -- CP-element group 459:  fork  transition  input  output  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	442 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459: 	468 
    -- CP-element group 459:  members (9) 
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_update_completed_
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_Update/$exit
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3034_Update/ca
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_sample_start_
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_Sample/$entry
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_Sample/rr
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_sample_start_
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_Sample/$entry
      -- CP-element group 459: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_Sample/rr
      -- 
    ca_7179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3034_inst_ack_1, ack => zeropad3D_CP_2067_elements(459)); -- 
    rr_7187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(459), ack => type_cast_3098_inst_req_0); -- 
    rr_7297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(459), ack => type_cast_3123_inst_req_0); -- 
    -- CP-element group 460:  transition  input  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_sample_completed_
      -- CP-element group 460: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_Sample/$exit
      -- CP-element group 460: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_Sample/ra
      -- 
    ra_7188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3098_inst_ack_0, ack => zeropad3D_CP_2067_elements(460)); -- 
    -- CP-element group 461:  transition  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	442 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (16) 
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_update_completed_
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_Update/$exit
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3098_Update/ca
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_resized_1
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_scaled_1
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_computed_1
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_resize_1/$entry
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_resize_1/$exit
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_resize_1/index_resize_req
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_resize_1/index_resize_ack
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_scale_1/$entry
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_scale_1/$exit
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_scale_1/scale_rename_req
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_index_scale_1/scale_rename_ack
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_Sample/req
      -- 
    ca_7193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3098_inst_ack_1, ack => zeropad3D_CP_2067_elements(461)); -- 
    req_7218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(461), ack => array_obj_ref_3104_index_offset_req_0); -- 
    -- CP-element group 462:  transition  input  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	477 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_sample_complete
      -- CP-element group 462: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_Sample/$exit
      -- CP-element group 462: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_Sample/ack
      -- 
    ack_7219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3104_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(462)); -- 
    -- CP-element group 463:  transition  input  output  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	442 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (11) 
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_root_address_calculated
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_offset_calculated
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_Update/$exit
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_final_index_sum_regn_Update/ack
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_base_plus_offset/$entry
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_base_plus_offset/$exit
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_base_plus_offset/sum_rename_req
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3104_base_plus_offset/sum_rename_ack
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_request/$entry
      -- CP-element group 463: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_request/req
      -- 
    ack_7224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3104_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(463)); -- 
    req_7233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(463), ack => addr_of_3105_final_reg_req_0); -- 
    -- CP-element group 464:  transition  input  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_request/$exit
      -- CP-element group 464: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_request/ack
      -- 
    ack_7234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3105_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(464)); -- 
    -- CP-element group 465:  join  fork  transition  input  output  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	442 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (24) 
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_complete/$exit
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3105_complete/ack
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_address_calculated
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_word_address_calculated
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_root_address_calculated
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_address_resized
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_addr_resize/$entry
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_addr_resize/$exit
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_addr_resize/base_resize_req
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_addr_resize/base_resize_ack
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_plus_offset/$entry
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_plus_offset/$exit
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_plus_offset/sum_rename_req
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_base_plus_offset/sum_rename_ack
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_word_addrgen/$entry
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_word_addrgen/$exit
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_word_addrgen/root_register_req
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_word_addrgen/root_register_ack
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Sample/word_access_start/$entry
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Sample/word_access_start/word_0/$entry
      -- CP-element group 465: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Sample/word_access_start/word_0/rr
      -- 
    ack_7239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3105_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(465)); -- 
    rr_7272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(465), ack => ptr_deref_3109_load_0_req_0); -- 
    -- CP-element group 466:  transition  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466:  members (5) 
      -- CP-element group 466: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_sample_completed_
      -- CP-element group 466: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Sample/$exit
      -- CP-element group 466: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Sample/word_access_start/$exit
      -- CP-element group 466: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Sample/word_access_start/word_0/$exit
      -- CP-element group 466: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Sample/word_access_start/word_0/ra
      -- 
    ra_7273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3109_load_0_ack_0, ack => zeropad3D_CP_2067_elements(466)); -- 
    -- CP-element group 467:  transition  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	442 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	474 
    -- CP-element group 467:  members (9) 
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_update_completed_
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/$exit
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/word_access_complete/$exit
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/word_access_complete/word_0/$exit
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/word_access_complete/word_0/ca
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/ptr_deref_3109_Merge/$entry
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/ptr_deref_3109_Merge/$exit
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/ptr_deref_3109_Merge/merge_req
      -- CP-element group 467: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3109_Update/ptr_deref_3109_Merge/merge_ack
      -- 
    ca_7284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3109_load_0_ack_1, ack => zeropad3D_CP_2067_elements(467)); -- 
    -- CP-element group 468:  transition  input  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	459 
    -- CP-element group 468: successors 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_sample_completed_
      -- CP-element group 468: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_Sample/$exit
      -- CP-element group 468: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_Sample/ra
      -- 
    ra_7298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3123_inst_ack_0, ack => zeropad3D_CP_2067_elements(468)); -- 
    -- CP-element group 469:  transition  input  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	442 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	470 
    -- CP-element group 469:  members (16) 
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_update_completed_
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_Update/$exit
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/type_cast_3123_Update/ca
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_resized_1
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_scaled_1
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_computed_1
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_resize_1/$entry
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_resize_1/$exit
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_resize_1/index_resize_req
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_resize_1/index_resize_ack
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_scale_1/$entry
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_scale_1/$exit
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_scale_1/scale_rename_req
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_index_scale_1/scale_rename_ack
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_Sample/req
      -- 
    ca_7303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3123_inst_ack_1, ack => zeropad3D_CP_2067_elements(469)); -- 
    req_7328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(469), ack => array_obj_ref_3129_index_offset_req_0); -- 
    -- CP-element group 470:  transition  input  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	469 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	477 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_sample_complete
      -- CP-element group 470: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_Sample/$exit
      -- CP-element group 470: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_Sample/ack
      -- 
    ack_7329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3129_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(470)); -- 
    -- CP-element group 471:  transition  input  output  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	442 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	472 
    -- CP-element group 471:  members (11) 
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_sample_start_
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_root_address_calculated
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_offset_calculated
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_Update/$exit
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_final_index_sum_regn_Update/ack
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_base_plus_offset/$entry
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_base_plus_offset/$exit
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_base_plus_offset/sum_rename_req
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/array_obj_ref_3129_base_plus_offset/sum_rename_ack
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_request/$entry
      -- CP-element group 471: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_request/req
      -- 
    ack_7334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3129_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(471)); -- 
    req_7343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(471), ack => addr_of_3130_final_reg_req_0); -- 
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	471 
    -- CP-element group 472: successors 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_sample_completed_
      -- CP-element group 472: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_request/$exit
      -- CP-element group 472: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_request/ack
      -- 
    ack_7344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3130_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(472)); -- 
    -- CP-element group 473:  fork  transition  input  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	442 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (19) 
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_update_completed_
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_complete/$exit
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/addr_of_3130_complete/ack
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_address_calculated
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_word_address_calculated
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_root_address_calculated
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_address_resized
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_addr_resize/$entry
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_addr_resize/$exit
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_addr_resize/base_resize_req
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_addr_resize/base_resize_ack
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_plus_offset/$entry
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_plus_offset/$exit
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_plus_offset/sum_rename_req
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_base_plus_offset/sum_rename_ack
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_word_addrgen/$entry
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_word_addrgen/$exit
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_word_addrgen/root_register_req
      -- CP-element group 473: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_word_addrgen/root_register_ack
      -- 
    ack_7349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3130_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(473)); -- 
    -- CP-element group 474:  join  transition  output  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	467 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (9) 
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_sample_start_
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/$entry
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/ptr_deref_3133_Split/$entry
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/ptr_deref_3133_Split/$exit
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/ptr_deref_3133_Split/split_req
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/ptr_deref_3133_Split/split_ack
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/word_access_start/$entry
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/word_access_start/word_0/$entry
      -- CP-element group 474: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/word_access_start/word_0/rr
      -- 
    rr_7387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(474), ack => ptr_deref_3133_store_0_req_0); -- 
    zeropad3D_cp_element_group_474: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_474"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(467) & zeropad3D_CP_2067_elements(473);
      gj_zeropad3D_cp_element_group_474 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(474), clk => clk, reset => reset); --
    end block;
    -- CP-element group 475:  transition  input  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475:  members (5) 
      -- CP-element group 475: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_sample_completed_
      -- CP-element group 475: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/$exit
      -- CP-element group 475: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/word_access_start/$exit
      -- CP-element group 475: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/word_access_start/word_0/$exit
      -- CP-element group 475: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Sample/word_access_start/word_0/ra
      -- 
    ra_7388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3133_store_0_ack_0, ack => zeropad3D_CP_2067_elements(475)); -- 
    -- CP-element group 476:  transition  input  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	442 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	477 
    -- CP-element group 476:  members (5) 
      -- CP-element group 476: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_update_completed_
      -- CP-element group 476: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Update/$exit
      -- CP-element group 476: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Update/word_access_complete/$exit
      -- CP-element group 476: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Update/word_access_complete/word_0/$exit
      -- CP-element group 476: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/ptr_deref_3133_Update/word_access_complete/word_0/ca
      -- 
    ca_7399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3133_store_0_ack_1, ack => zeropad3D_CP_2067_elements(476)); -- 
    -- CP-element group 477:  join  transition  place  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	462 
    -- CP-element group 477: 	470 
    -- CP-element group 477: 	476 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	1047 
    -- CP-element group 477:  members (5) 
      -- CP-element group 477: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135__exit__
      -- CP-element group 477: 	 branch_block_stmt_655/ifx_xelse946_ifx_xend994
      -- CP-element group 477: 	 branch_block_stmt_655/assign_stmt_3035_to_assign_stmt_3135/$exit
      -- CP-element group 477: 	 branch_block_stmt_655/ifx_xelse946_ifx_xend994_PhiReq/$entry
      -- CP-element group 477: 	 branch_block_stmt_655/ifx_xelse946_ifx_xend994_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_477: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_477"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(462) & zeropad3D_CP_2067_elements(470) & zeropad3D_CP_2067_elements(476);
      gj_zeropad3D_cp_element_group_477 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(477), clk => clk, reset => reset); --
    end block;
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	1047 
    -- CP-element group 478: successors 
    -- CP-element group 478:  members (3) 
      -- CP-element group 478: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_sample_completed_
      -- CP-element group 478: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_Sample/$exit
      -- CP-element group 478: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_Sample/ra
      -- 
    ra_7411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3141_inst_ack_0, ack => zeropad3D_CP_2067_elements(478)); -- 
    -- CP-element group 479:  branch  transition  place  input  output  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	1047 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479: 	481 
    -- CP-element group 479:  members (13) 
      -- CP-element group 479: 	 branch_block_stmt_655/if_stmt_3156__entry__
      -- CP-element group 479: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155__exit__
      -- CP-element group 479: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/$exit
      -- CP-element group 479: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_update_completed_
      -- CP-element group 479: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_Update/$exit
      -- CP-element group 479: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_Update/ca
      -- CP-element group 479: 	 branch_block_stmt_655/if_stmt_3156_dead_link/$entry
      -- CP-element group 479: 	 branch_block_stmt_655/if_stmt_3156_eval_test/$entry
      -- CP-element group 479: 	 branch_block_stmt_655/if_stmt_3156_eval_test/$exit
      -- CP-element group 479: 	 branch_block_stmt_655/if_stmt_3156_eval_test/branch_req
      -- CP-element group 479: 	 branch_block_stmt_655/R_cmp1002_3157_place
      -- CP-element group 479: 	 branch_block_stmt_655/if_stmt_3156_if_link/$entry
      -- CP-element group 479: 	 branch_block_stmt_655/if_stmt_3156_else_link/$entry
      -- 
    ca_7416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3141_inst_ack_1, ack => zeropad3D_CP_2067_elements(479)); -- 
    branch_req_7424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(479), ack => if_stmt_3156_branch_req_0); -- 
    -- CP-element group 480:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	1056 
    -- CP-element group 480: 	1057 
    -- CP-element group 480: 	1059 
    -- CP-element group 480: 	1060 
    -- CP-element group 480: 	1062 
    -- CP-element group 480: 	1063 
    -- CP-element group 480:  members (40) 
      -- CP-element group 480: 	 branch_block_stmt_655/merge_stmt_3162__exit__
      -- CP-element group 480: 	 branch_block_stmt_655/assign_stmt_3168__entry__
      -- CP-element group 480: 	 branch_block_stmt_655/assign_stmt_3168__exit__
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047
      -- CP-element group 480: 	 branch_block_stmt_655/if_stmt_3156_if_link/$exit
      -- CP-element group 480: 	 branch_block_stmt_655/if_stmt_3156_if_link/if_choice_transition
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xend994_ifx_xthen1004
      -- CP-element group 480: 	 branch_block_stmt_655/assign_stmt_3168/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/assign_stmt_3168/$exit
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xend994_ifx_xthen1004_PhiReq/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xend994_ifx_xthen1004_PhiReq/$exit
      -- CP-element group 480: 	 branch_block_stmt_655/merge_stmt_3162_PhiReqMerge
      -- CP-element group 480: 	 branch_block_stmt_655/merge_stmt_3162_PhiAck/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/merge_stmt_3162_PhiAck/$exit
      -- CP-element group 480: 	 branch_block_stmt_655/merge_stmt_3162_PhiAck/dummy
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/Sample/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/Sample/rr
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/Update/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/Update/cr
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/Sample/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/Sample/rr
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/Update/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/Update/cr
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/Sample/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/Sample/rr
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/Update/$entry
      -- CP-element group 480: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3156_branch_ack_1, ack => zeropad3D_CP_2067_elements(480)); -- 
    rr_12622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(480), ack => type_cast_3280_inst_req_0); -- 
    cr_12627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(480), ack => type_cast_3280_inst_req_1); -- 
    rr_12645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(480), ack => type_cast_3272_inst_req_0); -- 
    cr_12650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(480), ack => type_cast_3272_inst_req_1); -- 
    rr_12668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(480), ack => type_cast_3268_inst_req_0); -- 
    cr_12673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(480), ack => type_cast_3268_inst_req_1); -- 
    -- CP-element group 481:  fork  transition  place  input  output  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	479 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	482 
    -- CP-element group 481: 	483 
    -- CP-element group 481: 	484 
    -- CP-element group 481: 	485 
    -- CP-element group 481: 	487 
    -- CP-element group 481: 	490 
    -- CP-element group 481: 	492 
    -- CP-element group 481: 	493 
    -- CP-element group 481: 	494 
    -- CP-element group 481: 	496 
    -- CP-element group 481:  members (54) 
      -- CP-element group 481: 	 branch_block_stmt_655/merge_stmt_3170__exit__
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254__entry__
      -- CP-element group 481: 	 branch_block_stmt_655/if_stmt_3156_else_link/$exit
      -- CP-element group 481: 	 branch_block_stmt_655/if_stmt_3156_else_link/else_choice_transition
      -- CP-element group 481: 	 branch_block_stmt_655/ifx_xend994_ifx_xelse1009
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_sample_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_update_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_Sample/rr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_sample_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_update_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_word_address_calculated
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_root_address_calculated
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Sample/word_access_start/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Sample/word_access_start/word_0/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Sample/word_access_start/word_0/rr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/word_access_complete/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/word_access_complete/word_0/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/word_access_complete/word_0/cr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_update_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_update_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_update_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_sample_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_update_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_word_address_calculated
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_root_address_calculated
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Sample/word_access_start/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Sample/word_access_start/word_0/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Sample/word_access_start/word_0/rr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/word_access_complete/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/word_access_complete/word_0/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/word_access_complete/word_0/cr
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_update_start_
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_655/ifx_xend994_ifx_xelse1009_PhiReq/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/ifx_xend994_ifx_xelse1009_PhiReq/$exit
      -- CP-element group 481: 	 branch_block_stmt_655/merge_stmt_3170_PhiReqMerge
      -- CP-element group 481: 	 branch_block_stmt_655/merge_stmt_3170_PhiAck/$entry
      -- CP-element group 481: 	 branch_block_stmt_655/merge_stmt_3170_PhiAck/$exit
      -- CP-element group 481: 	 branch_block_stmt_655/merge_stmt_3170_PhiAck/dummy
      -- 
    else_choice_transition_7433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3156_branch_ack_0, ack => zeropad3D_CP_2067_elements(481)); -- 
    rr_7449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => type_cast_3180_inst_req_0); -- 
    cr_7454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => type_cast_3180_inst_req_1); -- 
    rr_7471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => LOAD_col_high_3183_load_0_req_0); -- 
    cr_7482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => LOAD_col_high_3183_load_0_req_1); -- 
    cr_7501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => type_cast_3187_inst_req_1); -- 
    cr_7515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => type_cast_3207_inst_req_1); -- 
    cr_7529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => type_cast_3224_inst_req_1); -- 
    rr_7546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => LOAD_row_high_3227_load_0_req_0); -- 
    cr_7557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => LOAD_row_high_3227_load_0_req_1); -- 
    cr_7576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(481), ack => type_cast_3231_inst_req_1); -- 
    -- CP-element group 482:  transition  input  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	481 
    -- CP-element group 482: successors 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_sample_completed_
      -- CP-element group 482: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_Sample/$exit
      -- CP-element group 482: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_Sample/ra
      -- 
    ra_7450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3180_inst_ack_0, ack => zeropad3D_CP_2067_elements(482)); -- 
    -- CP-element group 483:  transition  input  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	481 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	488 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_update_completed_
      -- CP-element group 483: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_Update/$exit
      -- CP-element group 483: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3180_Update/ca
      -- 
    ca_7455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3180_inst_ack_1, ack => zeropad3D_CP_2067_elements(483)); -- 
    -- CP-element group 484:  transition  input  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	481 
    -- CP-element group 484: successors 
    -- CP-element group 484:  members (5) 
      -- CP-element group 484: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_sample_completed_
      -- CP-element group 484: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Sample/word_access_start/$exit
      -- CP-element group 484: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Sample/word_access_start/word_0/$exit
      -- CP-element group 484: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Sample/word_access_start/word_0/ra
      -- 
    ra_7472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3183_load_0_ack_0, ack => zeropad3D_CP_2067_elements(484)); -- 
    -- CP-element group 485:  transition  input  output  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	481 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	486 
    -- CP-element group 485:  members (12) 
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_update_completed_
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/word_access_complete/$exit
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/word_access_complete/word_0/$exit
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/word_access_complete/word_0/ca
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/LOAD_col_high_3183_Merge/$entry
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/LOAD_col_high_3183_Merge/$exit
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/LOAD_col_high_3183_Merge/merge_req
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_col_high_3183_Update/LOAD_col_high_3183_Merge/merge_ack
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_sample_start_
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_Sample/$entry
      -- CP-element group 485: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_Sample/rr
      -- 
    ca_7483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3183_load_0_ack_1, ack => zeropad3D_CP_2067_elements(485)); -- 
    rr_7496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(485), ack => type_cast_3187_inst_req_0); -- 
    -- CP-element group 486:  transition  input  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	485 
    -- CP-element group 486: successors 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_sample_completed_
      -- CP-element group 486: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_Sample/$exit
      -- CP-element group 486: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_Sample/ra
      -- 
    ra_7497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3187_inst_ack_0, ack => zeropad3D_CP_2067_elements(486)); -- 
    -- CP-element group 487:  transition  input  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	481 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_update_completed_
      -- CP-element group 487: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_Update/$exit
      -- CP-element group 487: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3187_Update/ca
      -- 
    ca_7502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3187_inst_ack_1, ack => zeropad3D_CP_2067_elements(487)); -- 
    -- CP-element group 488:  join  transition  output  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	483 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_sample_start_
      -- CP-element group 488: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_Sample/$entry
      -- CP-element group 488: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_Sample/rr
      -- 
    rr_7510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(488), ack => type_cast_3207_inst_req_0); -- 
    zeropad3D_cp_element_group_488: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_488"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(483) & zeropad3D_CP_2067_elements(487);
      gj_zeropad3D_cp_element_group_488 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(488), clk => clk, reset => reset); --
    end block;
    -- CP-element group 489:  transition  input  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_sample_completed_
      -- CP-element group 489: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_Sample/$exit
      -- CP-element group 489: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_Sample/ra
      -- 
    ra_7511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3207_inst_ack_0, ack => zeropad3D_CP_2067_elements(489)); -- 
    -- CP-element group 490:  transition  input  output  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	481 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	491 
    -- CP-element group 490:  members (6) 
      -- CP-element group 490: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_update_completed_
      -- CP-element group 490: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_Update/$exit
      -- CP-element group 490: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3207_Update/ca
      -- CP-element group 490: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_sample_start_
      -- CP-element group 490: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_Sample/$entry
      -- CP-element group 490: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_Sample/rr
      -- 
    ca_7516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3207_inst_ack_1, ack => zeropad3D_CP_2067_elements(490)); -- 
    rr_7524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(490), ack => type_cast_3224_inst_req_0); -- 
    -- CP-element group 491:  transition  input  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	490 
    -- CP-element group 491: successors 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_sample_completed_
      -- CP-element group 491: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_Sample/ra
      -- 
    ra_7525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3224_inst_ack_0, ack => zeropad3D_CP_2067_elements(491)); -- 
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	481 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	497 
    -- CP-element group 492:  members (3) 
      -- CP-element group 492: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_update_completed_
      -- CP-element group 492: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3224_Update/ca
      -- 
    ca_7530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3224_inst_ack_1, ack => zeropad3D_CP_2067_elements(492)); -- 
    -- CP-element group 493:  transition  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	481 
    -- CP-element group 493: successors 
    -- CP-element group 493:  members (5) 
      -- CP-element group 493: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_sample_completed_
      -- CP-element group 493: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Sample/$exit
      -- CP-element group 493: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Sample/word_access_start/$exit
      -- CP-element group 493: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Sample/word_access_start/word_0/$exit
      -- CP-element group 493: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Sample/word_access_start/word_0/ra
      -- 
    ra_7547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3227_load_0_ack_0, ack => zeropad3D_CP_2067_elements(493)); -- 
    -- CP-element group 494:  transition  input  output  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	481 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (12) 
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_update_completed_
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/$exit
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/word_access_complete/$exit
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/word_access_complete/word_0/$exit
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/word_access_complete/word_0/ca
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/LOAD_row_high_3227_Merge/$entry
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/LOAD_row_high_3227_Merge/$exit
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/LOAD_row_high_3227_Merge/merge_req
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/LOAD_row_high_3227_Update/LOAD_row_high_3227_Merge/merge_ack
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_sample_start_
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_Sample/$entry
      -- CP-element group 494: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_Sample/rr
      -- 
    ca_7558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3227_load_0_ack_1, ack => zeropad3D_CP_2067_elements(494)); -- 
    rr_7571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(494), ack => type_cast_3231_inst_req_0); -- 
    -- CP-element group 495:  transition  input  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_sample_completed_
      -- CP-element group 495: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_Sample/$exit
      -- CP-element group 495: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_Sample/ra
      -- 
    ra_7572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3231_inst_ack_0, ack => zeropad3D_CP_2067_elements(495)); -- 
    -- CP-element group 496:  transition  input  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	481 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	497 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_update_completed_
      -- CP-element group 496: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_Update/$exit
      -- CP-element group 496: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/type_cast_3231_Update/ca
      -- 
    ca_7577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3231_inst_ack_1, ack => zeropad3D_CP_2067_elements(496)); -- 
    -- CP-element group 497:  branch  join  transition  place  output  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	492 
    -- CP-element group 497: 	496 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497: 	499 
    -- CP-element group 497:  members (10) 
      -- CP-element group 497: 	 branch_block_stmt_655/if_stmt_3255__entry__
      -- CP-element group 497: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254__exit__
      -- CP-element group 497: 	 branch_block_stmt_655/assign_stmt_3176_to_assign_stmt_3254/$exit
      -- CP-element group 497: 	 branch_block_stmt_655/if_stmt_3255_dead_link/$entry
      -- CP-element group 497: 	 branch_block_stmt_655/if_stmt_3255_eval_test/$entry
      -- CP-element group 497: 	 branch_block_stmt_655/if_stmt_3255_eval_test/$exit
      -- CP-element group 497: 	 branch_block_stmt_655/if_stmt_3255_eval_test/branch_req
      -- CP-element group 497: 	 branch_block_stmt_655/R_cmp1038_3256_place
      -- CP-element group 497: 	 branch_block_stmt_655/if_stmt_3255_if_link/$entry
      -- CP-element group 497: 	 branch_block_stmt_655/if_stmt_3255_else_link/$entry
      -- 
    branch_req_7585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(497), ack => if_stmt_3255_branch_req_0); -- 
    zeropad3D_cp_element_group_497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(492) & zeropad3D_CP_2067_elements(496);
      gj_zeropad3D_cp_element_group_497 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 498:  fork  transition  place  input  output  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	497 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	1071 
    -- CP-element group 498: 	1072 
    -- CP-element group 498: 	1074 
    -- CP-element group 498: 	1075 
    -- CP-element group 498: 	1077 
    -- CP-element group 498: 	1078 
    -- CP-element group 498:  members (28) 
      -- CP-element group 498: 	 branch_block_stmt_655/if_stmt_3255_if_link/$exit
      -- CP-element group 498: 	 branch_block_stmt_655/if_stmt_3255_if_link/if_choice_transition
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/Sample/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/Sample/rr
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/Update/cr
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/Sample/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/Sample/rr
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/Update/cr
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/Sample/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/Sample/rr
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3255_branch_ack_1, ack => zeropad3D_CP_2067_elements(498)); -- 
    rr_12701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(498), ack => type_cast_3295_inst_req_0); -- 
    cr_12706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(498), ack => type_cast_3295_inst_req_1); -- 
    rr_12724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(498), ack => type_cast_3291_inst_req_0); -- 
    cr_12729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(498), ack => type_cast_3291_inst_req_1); -- 
    rr_12747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(498), ack => type_cast_3287_inst_req_0); -- 
    cr_12752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(498), ack => type_cast_3287_inst_req_1); -- 
    -- CP-element group 499:  fork  transition  place  input  output  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	497 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	1048 
    -- CP-element group 499: 	1049 
    -- CP-element group 499: 	1051 
    -- CP-element group 499: 	1052 
    -- CP-element group 499: 	1054 
    -- CP-element group 499:  members (22) 
      -- CP-element group 499: 	 branch_block_stmt_655/if_stmt_3255_else_link/$exit
      -- CP-element group 499: 	 branch_block_stmt_655/if_stmt_3255_else_link/else_choice_transition
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/Sample/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/Sample/rr
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/Update/cr
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/Sample/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/Sample/rr
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/Update/cr
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3262/$entry
      -- CP-element group 499: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/$entry
      -- 
    else_choice_transition_7594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3255_branch_ack_0, ack => zeropad3D_CP_2067_elements(499)); -- 
    rr_12565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(499), ack => type_cast_3278_inst_req_0); -- 
    cr_12570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(499), ack => type_cast_3278_inst_req_1); -- 
    rr_12588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(499), ack => type_cast_3274_inst_req_0); -- 
    cr_12593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(499), ack => type_cast_3274_inst_req_1); -- 
    -- CP-element group 500:  transition  input  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	1084 
    -- CP-element group 500: successors 
    -- CP-element group 500:  members (3) 
      -- CP-element group 500: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_sample_completed_
      -- CP-element group 500: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_Sample/$exit
      -- CP-element group 500: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_Sample/ra
      -- 
    ra_7608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3299_inst_ack_0, ack => zeropad3D_CP_2067_elements(500)); -- 
    -- CP-element group 501:  transition  input  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	1084 
    -- CP-element group 501: successors 
    -- CP-element group 501: 	522 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_update_completed_
      -- CP-element group 501: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_Update/$exit
      -- CP-element group 501: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_Update/ca
      -- 
    ca_7613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3299_inst_ack_1, ack => zeropad3D_CP_2067_elements(501)); -- 
    -- CP-element group 502:  transition  input  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	1084 
    -- CP-element group 502: successors 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_sample_completed_
      -- CP-element group 502: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_Sample/$exit
      -- CP-element group 502: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_Sample/ra
      -- 
    ra_7622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3309_inst_ack_0, ack => zeropad3D_CP_2067_elements(502)); -- 
    -- CP-element group 503:  transition  input  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	1084 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	522 
    -- CP-element group 503:  members (3) 
      -- CP-element group 503: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_update_completed_
      -- CP-element group 503: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_Update/$exit
      -- CP-element group 503: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_Update/ca
      -- 
    ca_7627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3309_inst_ack_1, ack => zeropad3D_CP_2067_elements(503)); -- 
    -- CP-element group 504:  transition  input  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	1084 
    -- CP-element group 504: successors 
    -- CP-element group 504:  members (5) 
      -- CP-element group 504: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_sample_completed_
      -- CP-element group 504: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Sample/$exit
      -- CP-element group 504: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Sample/word_access_start/$exit
      -- CP-element group 504: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Sample/word_access_start/word_0/$exit
      -- CP-element group 504: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Sample/word_access_start/word_0/ra
      -- 
    ra_7644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3318_load_0_ack_0, ack => zeropad3D_CP_2067_elements(504)); -- 
    -- CP-element group 505:  transition  input  output  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	1084 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	518 
    -- CP-element group 505:  members (12) 
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_Sample/rr
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_Sample/$entry
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_sample_start_
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_update_completed_
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/$exit
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/word_access_complete/$exit
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/word_access_complete/word_0/$exit
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/word_access_complete/word_0/ca
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/LOAD_pad_3318_Merge/$entry
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/LOAD_pad_3318_Merge/$exit
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/LOAD_pad_3318_Merge/merge_req
      -- CP-element group 505: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/LOAD_pad_3318_Merge/merge_ack
      -- 
    ca_7655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3318_load_0_ack_1, ack => zeropad3D_CP_2067_elements(505)); -- 
    rr_7809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(505), ack => type_cast_3348_inst_req_0); -- 
    -- CP-element group 506:  transition  input  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	1084 
    -- CP-element group 506: successors 
    -- CP-element group 506:  members (5) 
      -- CP-element group 506: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_sample_completed_
      -- CP-element group 506: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Sample/$exit
      -- CP-element group 506: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Sample/word_access_start/$exit
      -- CP-element group 506: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Sample/word_access_start/word_0/$exit
      -- CP-element group 506: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Sample/word_access_start/word_0/ra
      -- 
    ra_7677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3321_load_0_ack_0, ack => zeropad3D_CP_2067_elements(506)); -- 
    -- CP-element group 507:  transition  input  output  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	1084 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	512 
    -- CP-element group 507:  members (12) 
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_update_completed_
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/$exit
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/word_access_complete/$exit
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/word_access_complete/word_0/$exit
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/word_access_complete/word_0/ca
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/LOAD_depth_high_3321_Merge/$entry
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/LOAD_depth_high_3321_Merge/$exit
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/LOAD_depth_high_3321_Merge/merge_req
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/LOAD_depth_high_3321_Merge/merge_ack
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_Sample/rr
      -- 
    ca_7688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3321_load_0_ack_1, ack => zeropad3D_CP_2067_elements(507)); -- 
    rr_7767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(507), ack => type_cast_3331_inst_req_0); -- 
    -- CP-element group 508:  transition  input  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	1084 
    -- CP-element group 508: successors 
    -- CP-element group 508:  members (5) 
      -- CP-element group 508: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_sample_completed_
      -- CP-element group 508: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Sample/$exit
      -- CP-element group 508: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Sample/word_access_start/$exit
      -- CP-element group 508: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Sample/word_access_start/word_0/$exit
      -- CP-element group 508: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Sample/word_access_start/word_0/ra
      -- 
    ra_7710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_3324_load_0_ack_0, ack => zeropad3D_CP_2067_elements(508)); -- 
    -- CP-element group 509:  fork  transition  input  output  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	1084 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	514 
    -- CP-element group 509: 	520 
    -- CP-element group 509:  members (15) 
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_Sample/$entry
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_sample_start_
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_Sample/rr
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_Sample/$entry
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_Sample/rr
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_sample_start_
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_update_completed_
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/$exit
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/word_access_complete/$exit
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/word_access_complete/word_0/$exit
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/word_access_complete/word_0/ca
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/LOAD_out_depth_high_3324_Merge/$entry
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/LOAD_out_depth_high_3324_Merge/$exit
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/LOAD_out_depth_high_3324_Merge/merge_req
      -- CP-element group 509: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/LOAD_out_depth_high_3324_Merge/merge_ack
      -- 
    ca_7721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_3324_load_0_ack_1, ack => zeropad3D_CP_2067_elements(509)); -- 
    rr_7781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(509), ack => type_cast_3335_inst_req_0); -- 
    rr_7823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(509), ack => type_cast_3352_inst_req_0); -- 
    -- CP-element group 510:  transition  input  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	1084 
    -- CP-element group 510: successors 
    -- CP-element group 510:  members (5) 
      -- CP-element group 510: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_sample_completed_
      -- CP-element group 510: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Sample/$exit
      -- CP-element group 510: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Sample/word_access_start/$exit
      -- CP-element group 510: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Sample/word_access_start/word_0/$exit
      -- CP-element group 510: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Sample/word_access_start/word_0/ra
      -- 
    ra_7743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_3327_load_0_ack_0, ack => zeropad3D_CP_2067_elements(510)); -- 
    -- CP-element group 511:  transition  input  output  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	1084 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	516 
    -- CP-element group 511:  members (12) 
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_Sample/rr
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_Sample/$entry
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_sample_start_
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_update_completed_
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/$exit
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/word_access_complete/$exit
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/word_access_complete/word_0/$exit
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/word_access_complete/word_0/ca
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/LOAD_out_col_high_3327_Merge/$entry
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/LOAD_out_col_high_3327_Merge/$exit
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/LOAD_out_col_high_3327_Merge/merge_req
      -- CP-element group 511: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/LOAD_out_col_high_3327_Merge/merge_ack
      -- 
    ca_7754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_3327_load_0_ack_1, ack => zeropad3D_CP_2067_elements(511)); -- 
    rr_7795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(511), ack => type_cast_3339_inst_req_0); -- 
    -- CP-element group 512:  transition  input  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	507 
    -- CP-element group 512: successors 
    -- CP-element group 512:  members (3) 
      -- CP-element group 512: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_sample_completed_
      -- CP-element group 512: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_Sample/$exit
      -- CP-element group 512: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_Sample/ra
      -- 
    ra_7768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 512_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3331_inst_ack_0, ack => zeropad3D_CP_2067_elements(512)); -- 
    -- CP-element group 513:  transition  input  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	1084 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	522 
    -- CP-element group 513:  members (3) 
      -- CP-element group 513: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_Update/ca
      -- CP-element group 513: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_Update/$exit
      -- CP-element group 513: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_update_completed_
      -- 
    ca_7773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3331_inst_ack_1, ack => zeropad3D_CP_2067_elements(513)); -- 
    -- CP-element group 514:  transition  input  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	509 
    -- CP-element group 514: successors 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_Sample/$exit
      -- CP-element group 514: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_sample_completed_
      -- CP-element group 514: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_Sample/ra
      -- 
    ra_7782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3335_inst_ack_0, ack => zeropad3D_CP_2067_elements(514)); -- 
    -- CP-element group 515:  transition  input  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	1084 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	522 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_update_completed_
      -- CP-element group 515: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_Update/ca
      -- CP-element group 515: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_Update/$exit
      -- 
    ca_7787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 515_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3335_inst_ack_1, ack => zeropad3D_CP_2067_elements(515)); -- 
    -- CP-element group 516:  transition  input  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	511 
    -- CP-element group 516: successors 
    -- CP-element group 516:  members (3) 
      -- CP-element group 516: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_Sample/ra
      -- CP-element group 516: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_Sample/$exit
      -- CP-element group 516: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_sample_completed_
      -- 
    ra_7796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3339_inst_ack_0, ack => zeropad3D_CP_2067_elements(516)); -- 
    -- CP-element group 517:  transition  input  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	1084 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	522 
    -- CP-element group 517:  members (3) 
      -- CP-element group 517: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_Update/ca
      -- CP-element group 517: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_Update/$exit
      -- CP-element group 517: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_update_completed_
      -- 
    ca_7801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3339_inst_ack_1, ack => zeropad3D_CP_2067_elements(517)); -- 
    -- CP-element group 518:  transition  input  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	505 
    -- CP-element group 518: successors 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_Sample/ra
      -- CP-element group 518: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_Sample/$exit
      -- CP-element group 518: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_sample_completed_
      -- 
    ra_7810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3348_inst_ack_0, ack => zeropad3D_CP_2067_elements(518)); -- 
    -- CP-element group 519:  transition  input  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	1084 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	522 
    -- CP-element group 519:  members (3) 
      -- CP-element group 519: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_Update/$exit
      -- CP-element group 519: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_Update/ca
      -- CP-element group 519: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_update_completed_
      -- 
    ca_7815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 519_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3348_inst_ack_1, ack => zeropad3D_CP_2067_elements(519)); -- 
    -- CP-element group 520:  transition  input  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	509 
    -- CP-element group 520: successors 
    -- CP-element group 520:  members (3) 
      -- CP-element group 520: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_Sample/ra
      -- CP-element group 520: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_Sample/$exit
      -- CP-element group 520: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_sample_completed_
      -- 
    ra_7824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3352_inst_ack_0, ack => zeropad3D_CP_2067_elements(520)); -- 
    -- CP-element group 521:  transition  input  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	1084 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	522 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_Update/ca
      -- CP-element group 521: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_Update/$exit
      -- CP-element group 521: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_update_completed_
      -- 
    ca_7829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3352_inst_ack_1, ack => zeropad3D_CP_2067_elements(521)); -- 
    -- CP-element group 522:  join  fork  transition  place  output  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	501 
    -- CP-element group 522: 	503 
    -- CP-element group 522: 	513 
    -- CP-element group 522: 	515 
    -- CP-element group 522: 	517 
    -- CP-element group 522: 	519 
    -- CP-element group 522: 	521 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	1095 
    -- CP-element group 522: 	1096 
    -- CP-element group 522: 	1097 
    -- CP-element group 522: 	1099 
    -- CP-element group 522: 	1100 
    -- CP-element group 522:  members (22) 
      -- CP-element group 522: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394__exit__
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/Sample/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/$exit
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/Update/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/Update/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/Update/cr
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3397/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/Sample/rr
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/Sample/rr
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/Sample/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/$entry
      -- CP-element group 522: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/Update/cr
      -- 
    cr_12865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(522), ack => type_cast_3409_inst_req_1); -- 
    rr_12860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(522), ack => type_cast_3409_inst_req_0); -- 
    rr_12883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(522), ack => type_cast_3413_inst_req_0); -- 
    cr_12888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(522), ack => type_cast_3413_inst_req_1); -- 
    zeropad3D_cp_element_group_522: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_522"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(501) & zeropad3D_CP_2067_elements(503) & zeropad3D_CP_2067_elements(513) & zeropad3D_CP_2067_elements(515) & zeropad3D_CP_2067_elements(517) & zeropad3D_CP_2067_elements(519) & zeropad3D_CP_2067_elements(521);
      gj_zeropad3D_cp_element_group_522 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(522), clk => clk, reset => reset); --
    end block;
    -- CP-element group 523:  transition  input  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	1107 
    -- CP-element group 523: successors 
    -- CP-element group 523:  members (3) 
      -- CP-element group 523: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_Sample/ra
      -- CP-element group 523: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_Sample/$exit
      -- CP-element group 523: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_sample_completed_
      -- 
    ra_7841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3420_inst_ack_0, ack => zeropad3D_CP_2067_elements(523)); -- 
    -- CP-element group 524:  branch  transition  place  input  output  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	1107 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	525 
    -- CP-element group 524: 	526 
    -- CP-element group 524:  members (13) 
      -- CP-element group 524: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428__exit__
      -- CP-element group 524: 	 branch_block_stmt_655/if_stmt_3429__entry__
      -- CP-element group 524: 	 branch_block_stmt_655/if_stmt_3429_else_link/$entry
      -- CP-element group 524: 	 branch_block_stmt_655/if_stmt_3429_if_link/$entry
      -- CP-element group 524: 	 branch_block_stmt_655/if_stmt_3429_eval_test/branch_req
      -- CP-element group 524: 	 branch_block_stmt_655/if_stmt_3429_eval_test/$exit
      -- CP-element group 524: 	 branch_block_stmt_655/if_stmt_3429_eval_test/$entry
      -- CP-element group 524: 	 branch_block_stmt_655/if_stmt_3429_dead_link/$entry
      -- CP-element group 524: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_Update/ca
      -- CP-element group 524: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_Update/$exit
      -- CP-element group 524: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_update_completed_
      -- CP-element group 524: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/$exit
      -- CP-element group 524: 	 branch_block_stmt_655/R_cmp1117_3430_place
      -- 
    ca_7846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3420_inst_ack_1, ack => zeropad3D_CP_2067_elements(524)); -- 
    branch_req_7854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(524), ack => if_stmt_3429_branch_req_0); -- 
    -- CP-element group 525:  transition  place  input  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	524 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	1108 
    -- CP-element group 525:  members (5) 
      -- CP-element group 525: 	 branch_block_stmt_655/if_stmt_3429_if_link/if_choice_transition
      -- CP-element group 525: 	 branch_block_stmt_655/if_stmt_3429_if_link/$exit
      -- CP-element group 525: 	 branch_block_stmt_655/whilex_xbody1112_ifx_xthen1148
      -- CP-element group 525: 	 branch_block_stmt_655/whilex_xbody1112_ifx_xthen1148_PhiReq/$entry
      -- CP-element group 525: 	 branch_block_stmt_655/whilex_xbody1112_ifx_xthen1148_PhiReq/$exit
      -- 
    if_choice_transition_7859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3429_branch_ack_1, ack => zeropad3D_CP_2067_elements(525)); -- 
    -- CP-element group 526:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	524 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	527 
    -- CP-element group 526: 	528 
    -- CP-element group 526: 	530 
    -- CP-element group 526:  members (27) 
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466__entry__
      -- CP-element group 526: 	 branch_block_stmt_655/merge_stmt_3435__exit__
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/word_access_complete/word_0/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/word_access_complete/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Sample/word_access_start/word_0/rr
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Sample/word_access_start/word_0/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Sample/word_access_start/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Sample/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_root_address_calculated
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_word_address_calculated
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_update_start_
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_sample_start_
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/if_stmt_3429_else_link/else_choice_transition
      -- CP-element group 526: 	 branch_block_stmt_655/if_stmt_3429_else_link/$exit
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_Update/cr
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_Update/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/whilex_xbody1112_lorx_xlhsx_xfalse1119
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_update_start_
      -- CP-element group 526: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/word_access_complete/word_0/cr
      -- CP-element group 526: 	 branch_block_stmt_655/merge_stmt_3435_PhiReqMerge
      -- CP-element group 526: 	 branch_block_stmt_655/merge_stmt_3435_PhiAck/dummy
      -- CP-element group 526: 	 branch_block_stmt_655/merge_stmt_3435_PhiAck/$exit
      -- CP-element group 526: 	 branch_block_stmt_655/merge_stmt_3435_PhiAck/$entry
      -- CP-element group 526: 	 branch_block_stmt_655/whilex_xbody1112_lorx_xlhsx_xfalse1119_PhiReq/$exit
      -- CP-element group 526: 	 branch_block_stmt_655/whilex_xbody1112_lorx_xlhsx_xfalse1119_PhiReq/$entry
      -- 
    else_choice_transition_7863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 526_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3429_branch_ack_0, ack => zeropad3D_CP_2067_elements(526)); -- 
    rr_7884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(526), ack => LOAD_row_high_3437_load_0_req_0); -- 
    cr_7914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(526), ack => type_cast_3441_inst_req_1); -- 
    cr_7895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(526), ack => LOAD_row_high_3437_load_0_req_1); -- 
    -- CP-element group 527:  transition  input  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	526 
    -- CP-element group 527: successors 
    -- CP-element group 527:  members (5) 
      -- CP-element group 527: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Sample/word_access_start/word_0/ra
      -- CP-element group 527: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Sample/word_access_start/word_0/$exit
      -- CP-element group 527: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Sample/word_access_start/$exit
      -- CP-element group 527: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Sample/$exit
      -- CP-element group 527: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_sample_completed_
      -- 
    ra_7885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3437_load_0_ack_0, ack => zeropad3D_CP_2067_elements(527)); -- 
    -- CP-element group 528:  transition  input  output  bypass 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	526 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	529 
    -- CP-element group 528:  members (12) 
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/word_access_complete/word_0/$exit
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/word_access_complete/$exit
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/$exit
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_update_completed_
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/LOAD_row_high_3437_Merge/merge_ack
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/LOAD_row_high_3437_Merge/merge_req
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/LOAD_row_high_3437_Merge/$exit
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/LOAD_row_high_3437_Merge/$entry
      -- CP-element group 528: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/LOAD_row_high_3437_Update/word_access_complete/word_0/ca
      -- 
    ca_7896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3437_load_0_ack_1, ack => zeropad3D_CP_2067_elements(528)); -- 
    rr_7909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(528), ack => type_cast_3441_inst_req_0); -- 
    -- CP-element group 529:  transition  input  bypass 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	528 
    -- CP-element group 529: successors 
    -- CP-element group 529:  members (3) 
      -- CP-element group 529: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_Sample/ra
      -- CP-element group 529: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_Sample/$exit
      -- CP-element group 529: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_sample_completed_
      -- 
    ra_7910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 529_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3441_inst_ack_0, ack => zeropad3D_CP_2067_elements(529)); -- 
    -- CP-element group 530:  branch  transition  place  input  output  bypass 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	526 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	531 
    -- CP-element group 530: 	532 
    -- CP-element group 530:  members (13) 
      -- CP-element group 530: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466__exit__
      -- CP-element group 530: 	 branch_block_stmt_655/if_stmt_3467__entry__
      -- CP-element group 530: 	 branch_block_stmt_655/if_stmt_3467_if_link/$entry
      -- CP-element group 530: 	 branch_block_stmt_655/if_stmt_3467_eval_test/branch_req
      -- CP-element group 530: 	 branch_block_stmt_655/if_stmt_3467_eval_test/$exit
      -- CP-element group 530: 	 branch_block_stmt_655/if_stmt_3467_eval_test/$entry
      -- CP-element group 530: 	 branch_block_stmt_655/if_stmt_3467_dead_link/$entry
      -- CP-element group 530: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/$exit
      -- CP-element group 530: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_Update/ca
      -- CP-element group 530: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_Update/$exit
      -- CP-element group 530: 	 branch_block_stmt_655/R_cmp1129_3468_place
      -- CP-element group 530: 	 branch_block_stmt_655/assign_stmt_3438_to_assign_stmt_3466/type_cast_3441_update_completed_
      -- CP-element group 530: 	 branch_block_stmt_655/if_stmt_3467_else_link/$entry
      -- 
    ca_7915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3441_inst_ack_1, ack => zeropad3D_CP_2067_elements(530)); -- 
    branch_req_7923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(530), ack => if_stmt_3467_branch_req_0); -- 
    -- CP-element group 531:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	530 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	533 
    -- CP-element group 531: 	534 
    -- CP-element group 531:  members (18) 
      -- CP-element group 531: 	 branch_block_stmt_655/merge_stmt_3473__exit__
      -- CP-element group 531: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485__entry__
      -- CP-element group 531: 	 branch_block_stmt_655/if_stmt_3467_if_link/if_choice_transition
      -- CP-element group 531: 	 branch_block_stmt_655/if_stmt_3467_if_link/$exit
      -- CP-element group 531: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1119_lorx_xlhsx_xfalse1131
      -- CP-element group 531: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_Update/cr
      -- CP-element group 531: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_Update/$entry
      -- CP-element group 531: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_Sample/rr
      -- CP-element group 531: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_Sample/$entry
      -- CP-element group 531: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_update_start_
      -- CP-element group 531: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_sample_start_
      -- CP-element group 531: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/$entry
      -- CP-element group 531: 	 branch_block_stmt_655/merge_stmt_3473_PhiReqMerge
      -- CP-element group 531: 	 branch_block_stmt_655/merge_stmt_3473_PhiAck/dummy
      -- CP-element group 531: 	 branch_block_stmt_655/merge_stmt_3473_PhiAck/$exit
      -- CP-element group 531: 	 branch_block_stmt_655/merge_stmt_3473_PhiAck/$entry
      -- CP-element group 531: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1119_lorx_xlhsx_xfalse1131_PhiReq/$exit
      -- CP-element group 531: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1119_lorx_xlhsx_xfalse1131_PhiReq/$entry
      -- 
    if_choice_transition_7928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3467_branch_ack_1, ack => zeropad3D_CP_2067_elements(531)); -- 
    cr_7950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(531), ack => type_cast_3477_inst_req_1); -- 
    rr_7945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(531), ack => type_cast_3477_inst_req_0); -- 
    -- CP-element group 532:  transition  place  input  bypass 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	530 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	1108 
    -- CP-element group 532:  members (5) 
      -- CP-element group 532: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1119_ifx_xthen1148
      -- CP-element group 532: 	 branch_block_stmt_655/if_stmt_3467_else_link/else_choice_transition
      -- CP-element group 532: 	 branch_block_stmt_655/if_stmt_3467_else_link/$exit
      -- CP-element group 532: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1119_ifx_xthen1148_PhiReq/$entry
      -- CP-element group 532: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1119_ifx_xthen1148_PhiReq/$exit
      -- 
    else_choice_transition_7932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 532_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3467_branch_ack_0, ack => zeropad3D_CP_2067_elements(532)); -- 
    -- CP-element group 533:  transition  input  bypass 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	531 
    -- CP-element group 533: successors 
    -- CP-element group 533:  members (3) 
      -- CP-element group 533: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_Sample/ra
      -- CP-element group 533: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_Sample/$exit
      -- CP-element group 533: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_sample_completed_
      -- 
    ra_7946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 533_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3477_inst_ack_0, ack => zeropad3D_CP_2067_elements(533)); -- 
    -- CP-element group 534:  branch  transition  place  input  output  bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	531 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	535 
    -- CP-element group 534: 	536 
    -- CP-element group 534:  members (13) 
      -- CP-element group 534: 	 branch_block_stmt_655/if_stmt_3486__entry__
      -- CP-element group 534: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485__exit__
      -- CP-element group 534: 	 branch_block_stmt_655/R_cmp1136_3487_place
      -- CP-element group 534: 	 branch_block_stmt_655/if_stmt_3486_else_link/$entry
      -- CP-element group 534: 	 branch_block_stmt_655/if_stmt_3486_if_link/$entry
      -- CP-element group 534: 	 branch_block_stmt_655/if_stmt_3486_eval_test/branch_req
      -- CP-element group 534: 	 branch_block_stmt_655/if_stmt_3486_eval_test/$exit
      -- CP-element group 534: 	 branch_block_stmt_655/if_stmt_3486_eval_test/$entry
      -- CP-element group 534: 	 branch_block_stmt_655/if_stmt_3486_dead_link/$entry
      -- CP-element group 534: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_Update/ca
      -- CP-element group 534: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_Update/$exit
      -- CP-element group 534: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/type_cast_3477_update_completed_
      -- CP-element group 534: 	 branch_block_stmt_655/assign_stmt_3478_to_assign_stmt_3485/$exit
      -- 
    ca_7951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3477_inst_ack_1, ack => zeropad3D_CP_2067_elements(534)); -- 
    branch_req_7959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(534), ack => if_stmt_3486_branch_req_0); -- 
    -- CP-element group 535:  transition  place  input  bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	534 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	1108 
    -- CP-element group 535:  members (5) 
      -- CP-element group 535: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1131_ifx_xthen1148
      -- CP-element group 535: 	 branch_block_stmt_655/if_stmt_3486_if_link/if_choice_transition
      -- CP-element group 535: 	 branch_block_stmt_655/if_stmt_3486_if_link/$exit
      -- CP-element group 535: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1131_ifx_xthen1148_PhiReq/$entry
      -- CP-element group 535: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1131_ifx_xthen1148_PhiReq/$exit
      -- 
    if_choice_transition_7964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 535_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3486_branch_ack_1, ack => zeropad3D_CP_2067_elements(535)); -- 
    -- CP-element group 536:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	534 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	537 
    -- CP-element group 536: 	538 
    -- CP-element group 536: 	540 
    -- CP-element group 536:  members (27) 
      -- CP-element group 536: 	 branch_block_stmt_655/merge_stmt_3492__exit__
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511__entry__
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Sample/word_access_start/word_0/rr
      -- CP-element group 536: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1131_lorx_xlhsx_xfalse1138
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Sample/word_access_start/word_0/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Sample/word_access_start/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Sample/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_root_address_calculated
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_word_address_calculated
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_update_start_
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_sample_start_
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/if_stmt_3486_else_link/else_choice_transition
      -- CP-element group 536: 	 branch_block_stmt_655/if_stmt_3486_else_link/$exit
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_update_start_
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/word_access_complete/word_0/cr
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/word_access_complete/word_0/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/word_access_complete/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1131_lorx_xlhsx_xfalse1138_PhiReq/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1131_lorx_xlhsx_xfalse1138_PhiReq/$exit
      -- CP-element group 536: 	 branch_block_stmt_655/merge_stmt_3492_PhiAck/$entry
      -- CP-element group 536: 	 branch_block_stmt_655/merge_stmt_3492_PhiAck/$exit
      -- CP-element group 536: 	 branch_block_stmt_655/merge_stmt_3492_PhiAck/dummy
      -- CP-element group 536: 	 branch_block_stmt_655/merge_stmt_3492_PhiReqMerge
      -- 
    else_choice_transition_7968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 536_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3486_branch_ack_0, ack => zeropad3D_CP_2067_elements(536)); -- 
    rr_7989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(536), ack => LOAD_col_high_3494_load_0_req_0); -- 
    cr_8019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(536), ack => type_cast_3498_inst_req_1); -- 
    cr_8000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(536), ack => LOAD_col_high_3494_load_0_req_1); -- 
    -- CP-element group 537:  transition  input  bypass 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	536 
    -- CP-element group 537: successors 
    -- CP-element group 537:  members (5) 
      -- CP-element group 537: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Sample/word_access_start/word_0/$exit
      -- CP-element group 537: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Sample/word_access_start/$exit
      -- CP-element group 537: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Sample/$exit
      -- CP-element group 537: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_sample_completed_
      -- CP-element group 537: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Sample/word_access_start/word_0/ra
      -- 
    ra_7990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3494_load_0_ack_0, ack => zeropad3D_CP_2067_elements(537)); -- 
    -- CP-element group 538:  transition  input  output  bypass 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	536 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	539 
    -- CP-element group 538:  members (12) 
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_update_completed_
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_Sample/rr
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_Sample/$entry
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_sample_start_
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/LOAD_col_high_3494_Merge/merge_ack
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/LOAD_col_high_3494_Merge/merge_req
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/LOAD_col_high_3494_Merge/$exit
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/LOAD_col_high_3494_Merge/$entry
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/word_access_complete/word_0/ca
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/word_access_complete/word_0/$exit
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/word_access_complete/$exit
      -- CP-element group 538: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/LOAD_col_high_3494_Update/$exit
      -- 
    ca_8001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 538_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3494_load_0_ack_1, ack => zeropad3D_CP_2067_elements(538)); -- 
    rr_8014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(538), ack => type_cast_3498_inst_req_0); -- 
    -- CP-element group 539:  transition  input  bypass 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	538 
    -- CP-element group 539: successors 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_Sample/ra
      -- CP-element group 539: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_Sample/$exit
      -- CP-element group 539: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_sample_completed_
      -- 
    ra_8015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 539_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3498_inst_ack_0, ack => zeropad3D_CP_2067_elements(539)); -- 
    -- CP-element group 540:  branch  transition  place  input  output  bypass 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	536 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	541 
    -- CP-element group 540: 	542 
    -- CP-element group 540:  members (13) 
      -- CP-element group 540: 	 branch_block_stmt_655/if_stmt_3512__entry__
      -- CP-element group 540: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511__exit__
      -- CP-element group 540: 	 branch_block_stmt_655/R_cmp1146_3513_place
      -- CP-element group 540: 	 branch_block_stmt_655/if_stmt_3512_else_link/$entry
      -- CP-element group 540: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/$exit
      -- CP-element group 540: 	 branch_block_stmt_655/if_stmt_3512_if_link/$entry
      -- CP-element group 540: 	 branch_block_stmt_655/if_stmt_3512_eval_test/branch_req
      -- CP-element group 540: 	 branch_block_stmt_655/if_stmt_3512_eval_test/$exit
      -- CP-element group 540: 	 branch_block_stmt_655/if_stmt_3512_eval_test/$entry
      -- CP-element group 540: 	 branch_block_stmt_655/if_stmt_3512_dead_link/$entry
      -- CP-element group 540: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_Update/ca
      -- CP-element group 540: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_Update/$exit
      -- CP-element group 540: 	 branch_block_stmt_655/assign_stmt_3495_to_assign_stmt_3511/type_cast_3498_update_completed_
      -- 
    ca_8020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3498_inst_ack_1, ack => zeropad3D_CP_2067_elements(540)); -- 
    branch_req_8028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(540), ack => if_stmt_3512_branch_req_0); -- 
    -- CP-element group 541:  fork  transition  place  input  output  bypass 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	540 
    -- CP-element group 541: successors 
    -- CP-element group 541: 	557 
    -- CP-element group 541: 	558 
    -- CP-element group 541: 	560 
    -- CP-element group 541: 	562 
    -- CP-element group 541: 	564 
    -- CP-element group 541: 	566 
    -- CP-element group 541: 	568 
    -- CP-element group 541: 	570 
    -- CP-element group 541: 	572 
    -- CP-element group 541: 	575 
    -- CP-element group 541:  members (46) 
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681__entry__
      -- CP-element group 541: 	 branch_block_stmt_655/merge_stmt_3576__exit__
      -- CP-element group 541: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1138_ifx_xelse1169
      -- CP-element group 541: 	 branch_block_stmt_655/if_stmt_3512_if_link/if_choice_transition
      -- CP-element group 541: 	 branch_block_stmt_655/if_stmt_3512_if_link/$exit
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_sample_start_
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_update_start_
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_Sample/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_Sample/rr
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_update_start_
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_update_start_
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_update_start
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_Update/req
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_complete/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_complete/req
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_update_start_
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/word_access_complete/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/word_access_complete/word_0/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/word_access_complete/word_0/cr
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_update_start_
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_Update/cr
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_update_start_
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_update_start
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_Update/req
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_complete/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_complete/req
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_update_start_
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Update/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Update/word_access_complete/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Update/word_access_complete/word_0/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Update/word_access_complete/word_0/cr
      -- CP-element group 541: 	 branch_block_stmt_655/merge_stmt_3576_PhiAck/dummy
      -- CP-element group 541: 	 branch_block_stmt_655/merge_stmt_3576_PhiAck/$exit
      -- CP-element group 541: 	 branch_block_stmt_655/merge_stmt_3576_PhiAck/$entry
      -- CP-element group 541: 	 branch_block_stmt_655/merge_stmt_3576_PhiReqMerge
      -- CP-element group 541: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1138_ifx_xelse1169_PhiReq/$exit
      -- CP-element group 541: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1138_ifx_xelse1169_PhiReq/$entry
      -- 
    if_choice_transition_8033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 541_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3512_branch_ack_1, ack => zeropad3D_CP_2067_elements(541)); -- 
    rr_8191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => type_cast_3580_inst_req_0); -- 
    cr_8196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => type_cast_3580_inst_req_1); -- 
    cr_8210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => type_cast_3644_inst_req_1); -- 
    req_8241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => array_obj_ref_3650_index_offset_req_1); -- 
    req_8256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => addr_of_3651_final_reg_req_1); -- 
    cr_8301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => ptr_deref_3655_load_0_req_1); -- 
    cr_8320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => type_cast_3669_inst_req_1); -- 
    req_8351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => array_obj_ref_3675_index_offset_req_1); -- 
    req_8366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => addr_of_3676_final_reg_req_1); -- 
    cr_8416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(541), ack => ptr_deref_3679_store_0_req_1); -- 
    -- CP-element group 542:  transition  place  input  bypass 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	540 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	1108 
    -- CP-element group 542:  members (5) 
      -- CP-element group 542: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1138_ifx_xthen1148
      -- CP-element group 542: 	 branch_block_stmt_655/if_stmt_3512_else_link/else_choice_transition
      -- CP-element group 542: 	 branch_block_stmt_655/if_stmt_3512_else_link/$exit
      -- CP-element group 542: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1138_ifx_xthen1148_PhiReq/$entry
      -- CP-element group 542: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1138_ifx_xthen1148_PhiReq/$exit
      -- 
    else_choice_transition_8037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 542_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3512_branch_ack_0, ack => zeropad3D_CP_2067_elements(542)); -- 
    -- CP-element group 543:  transition  input  bypass 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	1108 
    -- CP-element group 543: successors 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_Sample/ra
      -- CP-element group 543: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_Sample/$exit
      -- CP-element group 543: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_sample_completed_
      -- 
    ra_8051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 543_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3522_inst_ack_0, ack => zeropad3D_CP_2067_elements(543)); -- 
    -- CP-element group 544:  transition  input  bypass 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	1108 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	547 
    -- CP-element group 544:  members (3) 
      -- CP-element group 544: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_Update/ca
      -- CP-element group 544: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_Update/$exit
      -- CP-element group 544: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_update_completed_
      -- 
    ca_8056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 544_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3522_inst_ack_1, ack => zeropad3D_CP_2067_elements(544)); -- 
    -- CP-element group 545:  transition  input  bypass 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	1108 
    -- CP-element group 545: successors 
    -- CP-element group 545:  members (3) 
      -- CP-element group 545: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_Sample/ra
      -- CP-element group 545: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_Sample/$exit
      -- CP-element group 545: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_sample_completed_
      -- 
    ra_8065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 545_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3527_inst_ack_0, ack => zeropad3D_CP_2067_elements(545)); -- 
    -- CP-element group 546:  transition  input  bypass 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	1108 
    -- CP-element group 546: successors 
    -- CP-element group 546: 	547 
    -- CP-element group 546:  members (3) 
      -- CP-element group 546: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_Update/ca
      -- CP-element group 546: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_Update/$exit
      -- CP-element group 546: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_update_completed_
      -- 
    ca_8070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 546_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3527_inst_ack_1, ack => zeropad3D_CP_2067_elements(546)); -- 
    -- CP-element group 547:  join  transition  output  bypass 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	544 
    -- CP-element group 547: 	546 
    -- CP-element group 547: successors 
    -- CP-element group 547: 	548 
    -- CP-element group 547:  members (3) 
      -- CP-element group 547: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_Sample/rr
      -- CP-element group 547: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_Sample/$entry
      -- CP-element group 547: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_sample_start_
      -- 
    rr_8078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(547), ack => type_cast_3561_inst_req_0); -- 
    zeropad3D_cp_element_group_547: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_547"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(544) & zeropad3D_CP_2067_elements(546);
      gj_zeropad3D_cp_element_group_547 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(547), clk => clk, reset => reset); --
    end block;
    -- CP-element group 548:  transition  input  bypass 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	547 
    -- CP-element group 548: successors 
    -- CP-element group 548:  members (3) 
      -- CP-element group 548: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_Sample/ra
      -- CP-element group 548: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_Sample/$exit
      -- CP-element group 548: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_sample_completed_
      -- 
    ra_8079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 548_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3561_inst_ack_0, ack => zeropad3D_CP_2067_elements(548)); -- 
    -- CP-element group 549:  transition  input  output  bypass 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	1108 
    -- CP-element group 549: successors 
    -- CP-element group 549: 	550 
    -- CP-element group 549:  members (16) 
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_resize_1/index_resize_req
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_resize_1/$exit
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_resize_1/$entry
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_computed_1
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_scaled_1
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_resized_1
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_Sample/req
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_Sample/$entry
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_Update/ca
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_Update/$exit
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_scale_1/scale_rename_ack
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_scale_1/scale_rename_req
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_scale_1/$exit
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_update_completed_
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_scale_1/$entry
      -- CP-element group 549: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_index_resize_1/index_resize_ack
      -- 
    ca_8084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 549_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3561_inst_ack_1, ack => zeropad3D_CP_2067_elements(549)); -- 
    req_8109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(549), ack => array_obj_ref_3567_index_offset_req_0); -- 
    -- CP-element group 550:  transition  input  bypass 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	549 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	556 
    -- CP-element group 550:  members (3) 
      -- CP-element group 550: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_Sample/ack
      -- CP-element group 550: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_Sample/$exit
      -- CP-element group 550: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_sample_complete
      -- 
    ack_8110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 550_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3567_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(550)); -- 
    -- CP-element group 551:  transition  input  output  bypass 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	1108 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	552 
    -- CP-element group 551:  members (11) 
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_Update/$exit
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_offset_calculated
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_root_address_calculated
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_sample_start_
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_request/req
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_request/$entry
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_base_plus_offset/sum_rename_ack
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_base_plus_offset/sum_rename_req
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_base_plus_offset/$exit
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_base_plus_offset/$entry
      -- CP-element group 551: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_Update/ack
      -- 
    ack_8115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 551_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3567_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(551)); -- 
    req_8124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(551), ack => addr_of_3568_final_reg_req_0); -- 
    -- CP-element group 552:  transition  input  bypass 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	551 
    -- CP-element group 552: successors 
    -- CP-element group 552:  members (3) 
      -- CP-element group 552: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_sample_completed_
      -- CP-element group 552: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_request/ack
      -- CP-element group 552: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_request/$exit
      -- 
    ack_8125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3568_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(552)); -- 
    -- CP-element group 553:  join  fork  transition  input  output  bypass 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	1108 
    -- CP-element group 553: successors 
    -- CP-element group 553: 	554 
    -- CP-element group 553:  members (28) 
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_word_addrgen/$entry
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_addr_resize/$exit
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/word_access_start/word_0/$entry
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_addr_resize/$entry
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_address_resized
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_root_address_calculated
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_word_addrgen/$exit
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_word_address_calculated
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/word_access_start/$entry
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_address_calculated
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/ptr_deref_3571_Split/split_ack
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_update_completed_
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_plus_offset/sum_rename_ack
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/ptr_deref_3571_Split/split_req
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_sample_start_
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_complete/ack
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/ptr_deref_3571_Split/$exit
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_plus_offset/sum_rename_req
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_complete/$exit
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/ptr_deref_3571_Split/$entry
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/$entry
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_plus_offset/$exit
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_word_addrgen/root_register_ack
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_plus_offset/$entry
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_addr_resize/base_resize_ack
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_word_addrgen/root_register_req
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/word_access_start/word_0/rr
      -- CP-element group 553: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_base_addr_resize/base_resize_req
      -- 
    ack_8130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3568_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(553)); -- 
    rr_8168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(553), ack => ptr_deref_3571_store_0_req_0); -- 
    -- CP-element group 554:  transition  input  bypass 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	553 
    -- CP-element group 554: successors 
    -- CP-element group 554:  members (5) 
      -- CP-element group 554: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/word_access_start/$exit
      -- CP-element group 554: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_sample_completed_
      -- CP-element group 554: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/$exit
      -- CP-element group 554: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/word_access_start/word_0/$exit
      -- CP-element group 554: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Sample/word_access_start/word_0/ra
      -- 
    ra_8169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 554_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3571_store_0_ack_0, ack => zeropad3D_CP_2067_elements(554)); -- 
    -- CP-element group 555:  transition  input  bypass 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	1108 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	556 
    -- CP-element group 555:  members (5) 
      -- CP-element group 555: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_update_completed_
      -- CP-element group 555: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Update/$exit
      -- CP-element group 555: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Update/word_access_complete/$exit
      -- CP-element group 555: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Update/word_access_complete/word_0/$exit
      -- CP-element group 555: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Update/word_access_complete/word_0/ca
      -- 
    ca_8180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 555_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3571_store_0_ack_1, ack => zeropad3D_CP_2067_elements(555)); -- 
    -- CP-element group 556:  join  transition  place  bypass 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	550 
    -- CP-element group 556: 	555 
    -- CP-element group 556: successors 
    -- CP-element group 556: 	1109 
    -- CP-element group 556:  members (5) 
      -- CP-element group 556: 	 branch_block_stmt_655/ifx_xthen1148_ifx_xend1217
      -- CP-element group 556: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574__exit__
      -- CP-element group 556: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/$exit
      -- CP-element group 556: 	 branch_block_stmt_655/ifx_xthen1148_ifx_xend1217_PhiReq/$exit
      -- CP-element group 556: 	 branch_block_stmt_655/ifx_xthen1148_ifx_xend1217_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_556: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_556"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(550) & zeropad3D_CP_2067_elements(555);
      gj_zeropad3D_cp_element_group_556 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(556), clk => clk, reset => reset); --
    end block;
    -- CP-element group 557:  transition  input  bypass 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	541 
    -- CP-element group 557: successors 
    -- CP-element group 557:  members (3) 
      -- CP-element group 557: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_sample_completed_
      -- CP-element group 557: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_Sample/$exit
      -- CP-element group 557: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_Sample/ra
      -- 
    ra_8192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 557_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3580_inst_ack_0, ack => zeropad3D_CP_2067_elements(557)); -- 
    -- CP-element group 558:  fork  transition  input  output  bypass 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	541 
    -- CP-element group 558: successors 
    -- CP-element group 558: 	559 
    -- CP-element group 558: 	567 
    -- CP-element group 558:  members (9) 
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_update_completed_
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_Update/$exit
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3580_Update/ca
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_sample_start_
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_Sample/$entry
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_Sample/rr
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_sample_start_
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_Sample/$entry
      -- CP-element group 558: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_Sample/rr
      -- 
    ca_8197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 558_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3580_inst_ack_1, ack => zeropad3D_CP_2067_elements(558)); -- 
    rr_8205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(558), ack => type_cast_3644_inst_req_0); -- 
    rr_8315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(558), ack => type_cast_3669_inst_req_0); -- 
    -- CP-element group 559:  transition  input  bypass 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: 	558 
    -- CP-element group 559: successors 
    -- CP-element group 559:  members (3) 
      -- CP-element group 559: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_sample_completed_
      -- CP-element group 559: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_Sample/$exit
      -- CP-element group 559: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_Sample/ra
      -- 
    ra_8206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 559_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3644_inst_ack_0, ack => zeropad3D_CP_2067_elements(559)); -- 
    -- CP-element group 560:  transition  input  output  bypass 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	541 
    -- CP-element group 560: successors 
    -- CP-element group 560: 	561 
    -- CP-element group 560:  members (16) 
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_update_completed_
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_Update/$exit
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3644_Update/ca
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_resized_1
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_scaled_1
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_computed_1
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_resize_1/$entry
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_resize_1/$exit
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_resize_1/index_resize_req
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_resize_1/index_resize_ack
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_scale_1/$entry
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_scale_1/$exit
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_scale_1/scale_rename_req
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_index_scale_1/scale_rename_ack
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_Sample/$entry
      -- CP-element group 560: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_Sample/req
      -- 
    ca_8211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 560_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3644_inst_ack_1, ack => zeropad3D_CP_2067_elements(560)); -- 
    req_8236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(560), ack => array_obj_ref_3650_index_offset_req_0); -- 
    -- CP-element group 561:  transition  input  bypass 
    -- CP-element group 561: predecessors 
    -- CP-element group 561: 	560 
    -- CP-element group 561: successors 
    -- CP-element group 561: 	576 
    -- CP-element group 561:  members (3) 
      -- CP-element group 561: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_sample_complete
      -- CP-element group 561: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_Sample/$exit
      -- CP-element group 561: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_Sample/ack
      -- 
    ack_8237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 561_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3650_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(561)); -- 
    -- CP-element group 562:  transition  input  output  bypass 
    -- CP-element group 562: predecessors 
    -- CP-element group 562: 	541 
    -- CP-element group 562: successors 
    -- CP-element group 562: 	563 
    -- CP-element group 562:  members (11) 
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_root_address_calculated
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_offset_calculated
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_Update/$exit
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_final_index_sum_regn_Update/ack
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_base_plus_offset/$entry
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_base_plus_offset/$exit
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_base_plus_offset/sum_rename_req
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3650_base_plus_offset/sum_rename_ack
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_request/$entry
      -- CP-element group 562: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_request/req
      -- 
    ack_8242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 562_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3650_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(562)); -- 
    req_8251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(562), ack => addr_of_3651_final_reg_req_0); -- 
    -- CP-element group 563:  transition  input  bypass 
    -- CP-element group 563: predecessors 
    -- CP-element group 563: 	562 
    -- CP-element group 563: successors 
    -- CP-element group 563:  members (3) 
      -- CP-element group 563: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_sample_completed_
      -- CP-element group 563: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_request/$exit
      -- CP-element group 563: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_request/ack
      -- 
    ack_8252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 563_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3651_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(563)); -- 
    -- CP-element group 564:  join  fork  transition  input  output  bypass 
    -- CP-element group 564: predecessors 
    -- CP-element group 564: 	541 
    -- CP-element group 564: successors 
    -- CP-element group 564: 	565 
    -- CP-element group 564:  members (24) 
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_update_completed_
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_complete/$exit
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3651_complete/ack
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_sample_start_
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_address_calculated
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_word_address_calculated
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_root_address_calculated
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_address_resized
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_addr_resize/$entry
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_addr_resize/$exit
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_addr_resize/base_resize_req
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_addr_resize/base_resize_ack
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_plus_offset/$entry
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_plus_offset/$exit
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_plus_offset/sum_rename_req
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_base_plus_offset/sum_rename_ack
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_word_addrgen/$entry
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_word_addrgen/$exit
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_word_addrgen/root_register_req
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_word_addrgen/root_register_ack
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Sample/$entry
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Sample/word_access_start/$entry
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Sample/word_access_start/word_0/$entry
      -- CP-element group 564: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Sample/word_access_start/word_0/rr
      -- 
    ack_8257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 564_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3651_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(564)); -- 
    rr_8290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(564), ack => ptr_deref_3655_load_0_req_0); -- 
    -- CP-element group 565:  transition  input  bypass 
    -- CP-element group 565: predecessors 
    -- CP-element group 565: 	564 
    -- CP-element group 565: successors 
    -- CP-element group 565:  members (5) 
      -- CP-element group 565: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_sample_completed_
      -- CP-element group 565: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Sample/$exit
      -- CP-element group 565: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Sample/word_access_start/$exit
      -- CP-element group 565: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Sample/word_access_start/word_0/$exit
      -- CP-element group 565: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Sample/word_access_start/word_0/ra
      -- 
    ra_8291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 565_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3655_load_0_ack_0, ack => zeropad3D_CP_2067_elements(565)); -- 
    -- CP-element group 566:  transition  input  bypass 
    -- CP-element group 566: predecessors 
    -- CP-element group 566: 	541 
    -- CP-element group 566: successors 
    -- CP-element group 566: 	573 
    -- CP-element group 566:  members (9) 
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_update_completed_
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/$exit
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/word_access_complete/$exit
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/word_access_complete/word_0/$exit
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/word_access_complete/word_0/ca
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/ptr_deref_3655_Merge/$entry
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/ptr_deref_3655_Merge/$exit
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/ptr_deref_3655_Merge/merge_req
      -- CP-element group 566: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3655_Update/ptr_deref_3655_Merge/merge_ack
      -- 
    ca_8302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 566_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3655_load_0_ack_1, ack => zeropad3D_CP_2067_elements(566)); -- 
    -- CP-element group 567:  transition  input  bypass 
    -- CP-element group 567: predecessors 
    -- CP-element group 567: 	558 
    -- CP-element group 567: successors 
    -- CP-element group 567:  members (3) 
      -- CP-element group 567: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_sample_completed_
      -- CP-element group 567: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_Sample/$exit
      -- CP-element group 567: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_Sample/ra
      -- 
    ra_8316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 567_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3669_inst_ack_0, ack => zeropad3D_CP_2067_elements(567)); -- 
    -- CP-element group 568:  transition  input  output  bypass 
    -- CP-element group 568: predecessors 
    -- CP-element group 568: 	541 
    -- CP-element group 568: successors 
    -- CP-element group 568: 	569 
    -- CP-element group 568:  members (16) 
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_update_completed_
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_Update/$exit
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/type_cast_3669_Update/ca
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_resized_1
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_scaled_1
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_computed_1
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_resize_1/$entry
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_resize_1/$exit
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_resize_1/index_resize_req
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_resize_1/index_resize_ack
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_scale_1/$entry
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_scale_1/$exit
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_scale_1/scale_rename_req
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_index_scale_1/scale_rename_ack
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_Sample/$entry
      -- CP-element group 568: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_Sample/req
      -- 
    ca_8321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 568_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3669_inst_ack_1, ack => zeropad3D_CP_2067_elements(568)); -- 
    req_8346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(568), ack => array_obj_ref_3675_index_offset_req_0); -- 
    -- CP-element group 569:  transition  input  bypass 
    -- CP-element group 569: predecessors 
    -- CP-element group 569: 	568 
    -- CP-element group 569: successors 
    -- CP-element group 569: 	576 
    -- CP-element group 569:  members (3) 
      -- CP-element group 569: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_sample_complete
      -- CP-element group 569: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_Sample/$exit
      -- CP-element group 569: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_Sample/ack
      -- 
    ack_8347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 569_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3675_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(569)); -- 
    -- CP-element group 570:  transition  input  output  bypass 
    -- CP-element group 570: predecessors 
    -- CP-element group 570: 	541 
    -- CP-element group 570: successors 
    -- CP-element group 570: 	571 
    -- CP-element group 570:  members (11) 
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_sample_start_
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_root_address_calculated
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_offset_calculated
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_Update/$exit
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_final_index_sum_regn_Update/ack
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_base_plus_offset/$entry
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_base_plus_offset/$exit
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_base_plus_offset/sum_rename_req
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/array_obj_ref_3675_base_plus_offset/sum_rename_ack
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_request/$entry
      -- CP-element group 570: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_request/req
      -- 
    ack_8352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 570_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3675_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(570)); -- 
    req_8361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(570), ack => addr_of_3676_final_reg_req_0); -- 
    -- CP-element group 571:  transition  input  bypass 
    -- CP-element group 571: predecessors 
    -- CP-element group 571: 	570 
    -- CP-element group 571: successors 
    -- CP-element group 571:  members (3) 
      -- CP-element group 571: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_sample_completed_
      -- CP-element group 571: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_request/$exit
      -- CP-element group 571: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_request/ack
      -- 
    ack_8362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 571_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3676_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(571)); -- 
    -- CP-element group 572:  fork  transition  input  bypass 
    -- CP-element group 572: predecessors 
    -- CP-element group 572: 	541 
    -- CP-element group 572: successors 
    -- CP-element group 572: 	573 
    -- CP-element group 572:  members (19) 
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_update_completed_
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_complete/$exit
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/addr_of_3676_complete/ack
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_address_calculated
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_word_address_calculated
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_root_address_calculated
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_address_resized
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_addr_resize/$entry
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_addr_resize/$exit
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_addr_resize/base_resize_req
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_addr_resize/base_resize_ack
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_plus_offset/$entry
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_plus_offset/$exit
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_plus_offset/sum_rename_req
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_base_plus_offset/sum_rename_ack
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_word_addrgen/$entry
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_word_addrgen/$exit
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_word_addrgen/root_register_req
      -- CP-element group 572: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_word_addrgen/root_register_ack
      -- 
    ack_8367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 572_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3676_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(572)); -- 
    -- CP-element group 573:  join  transition  output  bypass 
    -- CP-element group 573: predecessors 
    -- CP-element group 573: 	566 
    -- CP-element group 573: 	572 
    -- CP-element group 573: successors 
    -- CP-element group 573: 	574 
    -- CP-element group 573:  members (9) 
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_sample_start_
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/$entry
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/ptr_deref_3679_Split/$entry
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/ptr_deref_3679_Split/$exit
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/ptr_deref_3679_Split/split_req
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/ptr_deref_3679_Split/split_ack
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/word_access_start/$entry
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/word_access_start/word_0/$entry
      -- CP-element group 573: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/word_access_start/word_0/rr
      -- 
    rr_8405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(573), ack => ptr_deref_3679_store_0_req_0); -- 
    zeropad3D_cp_element_group_573: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_573"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(566) & zeropad3D_CP_2067_elements(572);
      gj_zeropad3D_cp_element_group_573 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(573), clk => clk, reset => reset); --
    end block;
    -- CP-element group 574:  transition  input  bypass 
    -- CP-element group 574: predecessors 
    -- CP-element group 574: 	573 
    -- CP-element group 574: successors 
    -- CP-element group 574:  members (5) 
      -- CP-element group 574: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_sample_completed_
      -- CP-element group 574: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/$exit
      -- CP-element group 574: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/word_access_start/$exit
      -- CP-element group 574: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/word_access_start/word_0/$exit
      -- CP-element group 574: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Sample/word_access_start/word_0/ra
      -- 
    ra_8406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 574_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3679_store_0_ack_0, ack => zeropad3D_CP_2067_elements(574)); -- 
    -- CP-element group 575:  transition  input  bypass 
    -- CP-element group 575: predecessors 
    -- CP-element group 575: 	541 
    -- CP-element group 575: successors 
    -- CP-element group 575: 	576 
    -- CP-element group 575:  members (5) 
      -- CP-element group 575: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_update_completed_
      -- CP-element group 575: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Update/$exit
      -- CP-element group 575: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Update/word_access_complete/$exit
      -- CP-element group 575: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Update/word_access_complete/word_0/$exit
      -- CP-element group 575: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/ptr_deref_3679_Update/word_access_complete/word_0/ca
      -- 
    ca_8417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 575_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3679_store_0_ack_1, ack => zeropad3D_CP_2067_elements(575)); -- 
    -- CP-element group 576:  join  transition  place  bypass 
    -- CP-element group 576: predecessors 
    -- CP-element group 576: 	561 
    -- CP-element group 576: 	569 
    -- CP-element group 576: 	575 
    -- CP-element group 576: successors 
    -- CP-element group 576: 	1109 
    -- CP-element group 576:  members (5) 
      -- CP-element group 576: 	 branch_block_stmt_655/ifx_xelse1169_ifx_xend1217
      -- CP-element group 576: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681__exit__
      -- CP-element group 576: 	 branch_block_stmt_655/assign_stmt_3581_to_assign_stmt_3681/$exit
      -- CP-element group 576: 	 branch_block_stmt_655/ifx_xelse1169_ifx_xend1217_PhiReq/$entry
      -- CP-element group 576: 	 branch_block_stmt_655/ifx_xelse1169_ifx_xend1217_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_576: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_576"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(561) & zeropad3D_CP_2067_elements(569) & zeropad3D_CP_2067_elements(575);
      gj_zeropad3D_cp_element_group_576 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(576), clk => clk, reset => reset); --
    end block;
    -- CP-element group 577:  transition  input  bypass 
    -- CP-element group 577: predecessors 
    -- CP-element group 577: 	1109 
    -- CP-element group 577: successors 
    -- CP-element group 577:  members (3) 
      -- CP-element group 577: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_sample_completed_
      -- CP-element group 577: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_Sample/$exit
      -- CP-element group 577: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_Sample/ra
      -- 
    ra_8429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 577_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3687_inst_ack_0, ack => zeropad3D_CP_2067_elements(577)); -- 
    -- CP-element group 578:  branch  transition  place  input  output  bypass 
    -- CP-element group 578: predecessors 
    -- CP-element group 578: 	1109 
    -- CP-element group 578: successors 
    -- CP-element group 578: 	579 
    -- CP-element group 578: 	580 
    -- CP-element group 578:  members (13) 
      -- CP-element group 578: 	 branch_block_stmt_655/if_stmt_3702__entry__
      -- CP-element group 578: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701__exit__
      -- CP-element group 578: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/$exit
      -- CP-element group 578: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_update_completed_
      -- CP-element group 578: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_Update/$exit
      -- CP-element group 578: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_Update/ca
      -- CP-element group 578: 	 branch_block_stmt_655/if_stmt_3702_dead_link/$entry
      -- CP-element group 578: 	 branch_block_stmt_655/if_stmt_3702_eval_test/$entry
      -- CP-element group 578: 	 branch_block_stmt_655/if_stmt_3702_eval_test/$exit
      -- CP-element group 578: 	 branch_block_stmt_655/if_stmt_3702_eval_test/branch_req
      -- CP-element group 578: 	 branch_block_stmt_655/R_cmp1225_3703_place
      -- CP-element group 578: 	 branch_block_stmt_655/if_stmt_3702_if_link/$entry
      -- CP-element group 578: 	 branch_block_stmt_655/if_stmt_3702_else_link/$entry
      -- 
    ca_8434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 578_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3687_inst_ack_1, ack => zeropad3D_CP_2067_elements(578)); -- 
    branch_req_8442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(578), ack => if_stmt_3702_branch_req_0); -- 
    -- CP-element group 579:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 579: predecessors 
    -- CP-element group 579: 	578 
    -- CP-element group 579: successors 
    -- CP-element group 579: 	1118 
    -- CP-element group 579: 	1119 
    -- CP-element group 579: 	1121 
    -- CP-element group 579: 	1122 
    -- CP-element group 579: 	1124 
    -- CP-element group 579: 	1125 
    -- CP-element group 579:  members (40) 
      -- CP-element group 579: 	 branch_block_stmt_655/assign_stmt_3714__entry__
      -- CP-element group 579: 	 branch_block_stmt_655/merge_stmt_3708__exit__
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269
      -- CP-element group 579: 	 branch_block_stmt_655/assign_stmt_3714__exit__
      -- CP-element group 579: 	 branch_block_stmt_655/if_stmt_3702_if_link/$exit
      -- CP-element group 579: 	 branch_block_stmt_655/if_stmt_3702_if_link/if_choice_transition
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xend1217_ifx_xthen1227
      -- CP-element group 579: 	 branch_block_stmt_655/assign_stmt_3714/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/assign_stmt_3714/$exit
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/Sample/rr
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/Update/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/Sample/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/merge_stmt_3708_PhiAck/dummy
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/merge_stmt_3708_PhiAck/$exit
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/merge_stmt_3708_PhiAck/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/merge_stmt_3708_PhiReqMerge
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xend1217_ifx_xthen1227_PhiReq/$exit
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xend1217_ifx_xthen1227_PhiReq/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/Update/cr
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/Sample/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/Sample/rr
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/Update/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/Update/cr
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/Sample/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/Sample/rr
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/Update/$entry
      -- CP-element group 579: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/Update/cr
      -- 
    if_choice_transition_8447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 579_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3702_branch_ack_1, ack => zeropad3D_CP_2067_elements(579)); -- 
    rr_13073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(579), ack => type_cast_3804_inst_req_0); -- 
    cr_13078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(579), ack => type_cast_3804_inst_req_1); -- 
    rr_13096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(579), ack => type_cast_3811_inst_req_0); -- 
    cr_13101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(579), ack => type_cast_3811_inst_req_1); -- 
    rr_13119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(579), ack => type_cast_3817_inst_req_0); -- 
    cr_13124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(579), ack => type_cast_3817_inst_req_1); -- 
    -- CP-element group 580:  fork  transition  place  input  output  bypass 
    -- CP-element group 580: predecessors 
    -- CP-element group 580: 	578 
    -- CP-element group 580: successors 
    -- CP-element group 580: 	581 
    -- CP-element group 580: 	582 
    -- CP-element group 580: 	583 
    -- CP-element group 580: 	584 
    -- CP-element group 580: 	586 
    -- CP-element group 580: 	589 
    -- CP-element group 580: 	591 
    -- CP-element group 580: 	592 
    -- CP-element group 580: 	593 
    -- CP-element group 580: 	595 
    -- CP-element group 580:  members (54) 
      -- CP-element group 580: 	 branch_block_stmt_655/merge_stmt_3716__exit__
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793__entry__
      -- CP-element group 580: 	 branch_block_stmt_655/if_stmt_3702_else_link/$exit
      -- CP-element group 580: 	 branch_block_stmt_655/if_stmt_3702_else_link/else_choice_transition
      -- CP-element group 580: 	 branch_block_stmt_655/ifx_xend1217_ifx_xelse1232
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_sample_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_update_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_Sample/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_Sample/rr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_Update/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_Update/cr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_sample_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_update_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_word_address_calculated
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_root_address_calculated
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Sample/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Sample/word_access_start/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Sample/word_access_start/word_0/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Sample/word_access_start/word_0/rr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/word_access_complete/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/word_access_complete/word_0/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/word_access_complete/word_0/cr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_update_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_Update/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_Update/cr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_update_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_Update/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_Update/cr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_update_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_Update/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_Update/cr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_sample_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_update_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_word_address_calculated
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_root_address_calculated
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Sample/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Sample/word_access_start/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Sample/word_access_start/word_0/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Sample/word_access_start/word_0/rr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/word_access_complete/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/word_access_complete/word_0/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/word_access_complete/word_0/cr
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_update_start_
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_Update/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_Update/cr
      -- CP-element group 580: 	 branch_block_stmt_655/merge_stmt_3716_PhiAck/dummy
      -- CP-element group 580: 	 branch_block_stmt_655/merge_stmt_3716_PhiAck/$exit
      -- CP-element group 580: 	 branch_block_stmt_655/merge_stmt_3716_PhiAck/$entry
      -- CP-element group 580: 	 branch_block_stmt_655/merge_stmt_3716_PhiReqMerge
      -- CP-element group 580: 	 branch_block_stmt_655/ifx_xend1217_ifx_xelse1232_PhiReq/$exit
      -- CP-element group 580: 	 branch_block_stmt_655/ifx_xend1217_ifx_xelse1232_PhiReq/$entry
      -- 
    else_choice_transition_8451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 580_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3702_branch_ack_0, ack => zeropad3D_CP_2067_elements(580)); -- 
    rr_8467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => type_cast_3726_inst_req_0); -- 
    cr_8472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => type_cast_3726_inst_req_1); -- 
    rr_8489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => LOAD_col_high_3729_load_0_req_0); -- 
    cr_8500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => LOAD_col_high_3729_load_0_req_1); -- 
    cr_8519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => type_cast_3733_inst_req_1); -- 
    cr_8533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => type_cast_3747_inst_req_1); -- 
    cr_8547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => type_cast_3763_inst_req_1); -- 
    rr_8564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => LOAD_row_high_3766_load_0_req_0); -- 
    cr_8575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => LOAD_row_high_3766_load_0_req_1); -- 
    cr_8594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(580), ack => type_cast_3770_inst_req_1); -- 
    -- CP-element group 581:  transition  input  bypass 
    -- CP-element group 581: predecessors 
    -- CP-element group 581: 	580 
    -- CP-element group 581: successors 
    -- CP-element group 581:  members (3) 
      -- CP-element group 581: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_sample_completed_
      -- CP-element group 581: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_Sample/$exit
      -- CP-element group 581: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_Sample/ra
      -- 
    ra_8468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 581_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3726_inst_ack_0, ack => zeropad3D_CP_2067_elements(581)); -- 
    -- CP-element group 582:  transition  input  bypass 
    -- CP-element group 582: predecessors 
    -- CP-element group 582: 	580 
    -- CP-element group 582: successors 
    -- CP-element group 582: 	587 
    -- CP-element group 582:  members (3) 
      -- CP-element group 582: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_update_completed_
      -- CP-element group 582: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_Update/$exit
      -- CP-element group 582: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3726_Update/ca
      -- 
    ca_8473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 582_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3726_inst_ack_1, ack => zeropad3D_CP_2067_elements(582)); -- 
    -- CP-element group 583:  transition  input  bypass 
    -- CP-element group 583: predecessors 
    -- CP-element group 583: 	580 
    -- CP-element group 583: successors 
    -- CP-element group 583:  members (5) 
      -- CP-element group 583: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_sample_completed_
      -- CP-element group 583: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Sample/$exit
      -- CP-element group 583: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Sample/word_access_start/$exit
      -- CP-element group 583: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Sample/word_access_start/word_0/$exit
      -- CP-element group 583: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Sample/word_access_start/word_0/ra
      -- 
    ra_8490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 583_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3729_load_0_ack_0, ack => zeropad3D_CP_2067_elements(583)); -- 
    -- CP-element group 584:  transition  input  output  bypass 
    -- CP-element group 584: predecessors 
    -- CP-element group 584: 	580 
    -- CP-element group 584: successors 
    -- CP-element group 584: 	585 
    -- CP-element group 584:  members (12) 
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_update_completed_
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/$exit
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/word_access_complete/$exit
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/word_access_complete/word_0/$exit
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/word_access_complete/word_0/ca
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/LOAD_col_high_3729_Merge/$entry
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/LOAD_col_high_3729_Merge/$exit
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/LOAD_col_high_3729_Merge/merge_req
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_col_high_3729_Update/LOAD_col_high_3729_Merge/merge_ack
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_Sample/rr
      -- 
    ca_8501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 584_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3729_load_0_ack_1, ack => zeropad3D_CP_2067_elements(584)); -- 
    rr_8514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(584), ack => type_cast_3733_inst_req_0); -- 
    -- CP-element group 585:  transition  input  bypass 
    -- CP-element group 585: predecessors 
    -- CP-element group 585: 	584 
    -- CP-element group 585: successors 
    -- CP-element group 585:  members (3) 
      -- CP-element group 585: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_sample_completed_
      -- CP-element group 585: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_Sample/$exit
      -- CP-element group 585: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_Sample/ra
      -- 
    ra_8515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 585_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3733_inst_ack_0, ack => zeropad3D_CP_2067_elements(585)); -- 
    -- CP-element group 586:  transition  input  bypass 
    -- CP-element group 586: predecessors 
    -- CP-element group 586: 	580 
    -- CP-element group 586: successors 
    -- CP-element group 586: 	587 
    -- CP-element group 586:  members (3) 
      -- CP-element group 586: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_update_completed_
      -- CP-element group 586: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_Update/$exit
      -- CP-element group 586: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3733_Update/ca
      -- 
    ca_8520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 586_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3733_inst_ack_1, ack => zeropad3D_CP_2067_elements(586)); -- 
    -- CP-element group 587:  join  transition  output  bypass 
    -- CP-element group 587: predecessors 
    -- CP-element group 587: 	582 
    -- CP-element group 587: 	586 
    -- CP-element group 587: successors 
    -- CP-element group 587: 	588 
    -- CP-element group 587:  members (3) 
      -- CP-element group 587: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_sample_start_
      -- CP-element group 587: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_Sample/$entry
      -- CP-element group 587: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_Sample/rr
      -- 
    rr_8528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(587), ack => type_cast_3747_inst_req_0); -- 
    zeropad3D_cp_element_group_587: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_587"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(582) & zeropad3D_CP_2067_elements(586);
      gj_zeropad3D_cp_element_group_587 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(587), clk => clk, reset => reset); --
    end block;
    -- CP-element group 588:  transition  input  bypass 
    -- CP-element group 588: predecessors 
    -- CP-element group 588: 	587 
    -- CP-element group 588: successors 
    -- CP-element group 588:  members (3) 
      -- CP-element group 588: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_sample_completed_
      -- CP-element group 588: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_Sample/$exit
      -- CP-element group 588: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_Sample/ra
      -- 
    ra_8529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 588_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3747_inst_ack_0, ack => zeropad3D_CP_2067_elements(588)); -- 
    -- CP-element group 589:  transition  input  output  bypass 
    -- CP-element group 589: predecessors 
    -- CP-element group 589: 	580 
    -- CP-element group 589: successors 
    -- CP-element group 589: 	590 
    -- CP-element group 589:  members (6) 
      -- CP-element group 589: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_update_completed_
      -- CP-element group 589: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_Update/$exit
      -- CP-element group 589: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3747_Update/ca
      -- CP-element group 589: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_sample_start_
      -- CP-element group 589: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_Sample/$entry
      -- CP-element group 589: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_Sample/rr
      -- 
    ca_8534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 589_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3747_inst_ack_1, ack => zeropad3D_CP_2067_elements(589)); -- 
    rr_8542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(589), ack => type_cast_3763_inst_req_0); -- 
    -- CP-element group 590:  transition  input  bypass 
    -- CP-element group 590: predecessors 
    -- CP-element group 590: 	589 
    -- CP-element group 590: successors 
    -- CP-element group 590:  members (3) 
      -- CP-element group 590: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_sample_completed_
      -- CP-element group 590: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_Sample/$exit
      -- CP-element group 590: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_Sample/ra
      -- 
    ra_8543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 590_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3763_inst_ack_0, ack => zeropad3D_CP_2067_elements(590)); -- 
    -- CP-element group 591:  transition  input  bypass 
    -- CP-element group 591: predecessors 
    -- CP-element group 591: 	580 
    -- CP-element group 591: successors 
    -- CP-element group 591: 	596 
    -- CP-element group 591:  members (3) 
      -- CP-element group 591: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_update_completed_
      -- CP-element group 591: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_Update/$exit
      -- CP-element group 591: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3763_Update/ca
      -- 
    ca_8548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 591_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3763_inst_ack_1, ack => zeropad3D_CP_2067_elements(591)); -- 
    -- CP-element group 592:  transition  input  bypass 
    -- CP-element group 592: predecessors 
    -- CP-element group 592: 	580 
    -- CP-element group 592: successors 
    -- CP-element group 592:  members (5) 
      -- CP-element group 592: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_sample_completed_
      -- CP-element group 592: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Sample/$exit
      -- CP-element group 592: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Sample/word_access_start/$exit
      -- CP-element group 592: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Sample/word_access_start/word_0/$exit
      -- CP-element group 592: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Sample/word_access_start/word_0/ra
      -- 
    ra_8565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 592_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3766_load_0_ack_0, ack => zeropad3D_CP_2067_elements(592)); -- 
    -- CP-element group 593:  transition  input  output  bypass 
    -- CP-element group 593: predecessors 
    -- CP-element group 593: 	580 
    -- CP-element group 593: successors 
    -- CP-element group 593: 	594 
    -- CP-element group 593:  members (12) 
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_update_completed_
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/$exit
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/word_access_complete/$exit
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/word_access_complete/word_0/$exit
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/word_access_complete/word_0/ca
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/LOAD_row_high_3766_Merge/$entry
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/LOAD_row_high_3766_Merge/$exit
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/LOAD_row_high_3766_Merge/merge_req
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/LOAD_row_high_3766_Update/LOAD_row_high_3766_Merge/merge_ack
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_sample_start_
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_Sample/$entry
      -- CP-element group 593: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_Sample/rr
      -- 
    ca_8576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 593_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3766_load_0_ack_1, ack => zeropad3D_CP_2067_elements(593)); -- 
    rr_8589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(593), ack => type_cast_3770_inst_req_0); -- 
    -- CP-element group 594:  transition  input  bypass 
    -- CP-element group 594: predecessors 
    -- CP-element group 594: 	593 
    -- CP-element group 594: successors 
    -- CP-element group 594:  members (3) 
      -- CP-element group 594: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_sample_completed_
      -- CP-element group 594: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_Sample/$exit
      -- CP-element group 594: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_Sample/ra
      -- 
    ra_8590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 594_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3770_inst_ack_0, ack => zeropad3D_CP_2067_elements(594)); -- 
    -- CP-element group 595:  transition  input  bypass 
    -- CP-element group 595: predecessors 
    -- CP-element group 595: 	580 
    -- CP-element group 595: successors 
    -- CP-element group 595: 	596 
    -- CP-element group 595:  members (3) 
      -- CP-element group 595: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_update_completed_
      -- CP-element group 595: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_Update/$exit
      -- CP-element group 595: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/type_cast_3770_Update/ca
      -- 
    ca_8595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 595_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3770_inst_ack_1, ack => zeropad3D_CP_2067_elements(595)); -- 
    -- CP-element group 596:  branch  join  transition  place  output  bypass 
    -- CP-element group 596: predecessors 
    -- CP-element group 596: 	591 
    -- CP-element group 596: 	595 
    -- CP-element group 596: successors 
    -- CP-element group 596: 	597 
    -- CP-element group 596: 	598 
    -- CP-element group 596:  members (10) 
      -- CP-element group 596: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793__exit__
      -- CP-element group 596: 	 branch_block_stmt_655/if_stmt_3794__entry__
      -- CP-element group 596: 	 branch_block_stmt_655/assign_stmt_3722_to_assign_stmt_3793/$exit
      -- CP-element group 596: 	 branch_block_stmt_655/if_stmt_3794_dead_link/$entry
      -- CP-element group 596: 	 branch_block_stmt_655/if_stmt_3794_eval_test/$entry
      -- CP-element group 596: 	 branch_block_stmt_655/if_stmt_3794_eval_test/$exit
      -- CP-element group 596: 	 branch_block_stmt_655/if_stmt_3794_eval_test/branch_req
      -- CP-element group 596: 	 branch_block_stmt_655/R_cmp1260_3795_place
      -- CP-element group 596: 	 branch_block_stmt_655/if_stmt_3794_if_link/$entry
      -- CP-element group 596: 	 branch_block_stmt_655/if_stmt_3794_else_link/$entry
      -- 
    branch_req_8603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(596), ack => if_stmt_3794_branch_req_0); -- 
    zeropad3D_cp_element_group_596: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_596"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(591) & zeropad3D_CP_2067_elements(595);
      gj_zeropad3D_cp_element_group_596 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(596), clk => clk, reset => reset); --
    end block;
    -- CP-element group 597:  fork  transition  place  input  output  bypass 
    -- CP-element group 597: predecessors 
    -- CP-element group 597: 	596 
    -- CP-element group 597: successors 
    -- CP-element group 597: 	1133 
    -- CP-element group 597: 	1134 
    -- CP-element group 597: 	1136 
    -- CP-element group 597: 	1137 
    -- CP-element group 597:  members (20) 
      -- CP-element group 597: 	 branch_block_stmt_655/if_stmt_3794_if_link/$exit
      -- CP-element group 597: 	 branch_block_stmt_655/if_stmt_3794_if_link/if_choice_transition
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/Sample/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/Sample/rr
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/Update/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/Update/cr
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/Sample/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/Sample/rr
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/Update/$entry
      -- CP-element group 597: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/Update/cr
      -- 
    if_choice_transition_8608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 597_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3794_branch_ack_1, ack => zeropad3D_CP_2067_elements(597)); -- 
    rr_13152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(597), ack => type_cast_3826_inst_req_0); -- 
    cr_13157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(597), ack => type_cast_3826_inst_req_1); -- 
    rr_13175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(597), ack => type_cast_3830_inst_req_0); -- 
    cr_13180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(597), ack => type_cast_3830_inst_req_1); -- 
    -- CP-element group 598:  fork  transition  place  input  output  bypass 
    -- CP-element group 598: predecessors 
    -- CP-element group 598: 	596 
    -- CP-element group 598: successors 
    -- CP-element group 598: 	1110 
    -- CP-element group 598: 	1111 
    -- CP-element group 598: 	1112 
    -- CP-element group 598: 	1114 
    -- CP-element group 598: 	1115 
    -- CP-element group 598:  members (22) 
      -- CP-element group 598: 	 branch_block_stmt_655/if_stmt_3794_else_link/$exit
      -- CP-element group 598: 	 branch_block_stmt_655/if_stmt_3794_else_link/else_choice_transition
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/Sample/rr
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/Update/cr
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/Update/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3801/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/Sample/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/Update/cr
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/Update/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/Sample/rr
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/Sample/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/$entry
      -- CP-element group 598: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/$entry
      -- 
    else_choice_transition_8612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 598_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3794_branch_ack_0, ack => zeropad3D_CP_2067_elements(598)); -- 
    rr_13024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(598), ack => type_cast_3813_inst_req_0); -- 
    cr_13029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(598), ack => type_cast_3813_inst_req_1); -- 
    cr_13052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(598), ack => type_cast_3819_inst_req_1); -- 
    rr_13047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(598), ack => type_cast_3819_inst_req_0); -- 
    -- CP-element group 599:  transition  input  bypass 
    -- CP-element group 599: predecessors 
    -- CP-element group 599: 	1142 
    -- CP-element group 599: successors 
    -- CP-element group 599:  members (3) 
      -- CP-element group 599: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_sample_completed_
      -- CP-element group 599: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_Sample/$exit
      -- CP-element group 599: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_Sample/ra
      -- 
    ra_8626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 599_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3834_inst_ack_0, ack => zeropad3D_CP_2067_elements(599)); -- 
    -- CP-element group 600:  transition  input  bypass 
    -- CP-element group 600: predecessors 
    -- CP-element group 600: 	1142 
    -- CP-element group 600: successors 
    -- CP-element group 600: 	619 
    -- CP-element group 600:  members (3) 
      -- CP-element group 600: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_update_completed_
      -- CP-element group 600: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_Update/$exit
      -- CP-element group 600: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_Update/ca
      -- 
    ca_8631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 600_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3834_inst_ack_1, ack => zeropad3D_CP_2067_elements(600)); -- 
    -- CP-element group 601:  transition  input  bypass 
    -- CP-element group 601: predecessors 
    -- CP-element group 601: 	1142 
    -- CP-element group 601: successors 
    -- CP-element group 601:  members (5) 
      -- CP-element group 601: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_sample_completed_
      -- CP-element group 601: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Sample/$exit
      -- CP-element group 601: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Sample/word_access_start/$exit
      -- CP-element group 601: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Sample/word_access_start/word_0/$exit
      -- CP-element group 601: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Sample/word_access_start/word_0/ra
      -- 
    ra_8648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 601_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3849_load_0_ack_0, ack => zeropad3D_CP_2067_elements(601)); -- 
    -- CP-element group 602:  transition  input  output  bypass 
    -- CP-element group 602: predecessors 
    -- CP-element group 602: 	1142 
    -- CP-element group 602: successors 
    -- CP-element group 602: 	615 
    -- CP-element group 602:  members (12) 
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_update_completed_
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/$exit
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/word_access_complete/$exit
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/word_access_complete/word_0/$exit
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/word_access_complete/word_0/ca
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/LOAD_pad_3849_Merge/$entry
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/LOAD_pad_3849_Merge/$exit
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/LOAD_pad_3849_Merge/merge_req
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/LOAD_pad_3849_Merge/merge_ack
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_sample_start_
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_Sample/$entry
      -- CP-element group 602: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_Sample/rr
      -- 
    ca_8659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 602_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3849_load_0_ack_1, ack => zeropad3D_CP_2067_elements(602)); -- 
    rr_8813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(602), ack => type_cast_3879_inst_req_0); -- 
    -- CP-element group 603:  transition  input  bypass 
    -- CP-element group 603: predecessors 
    -- CP-element group 603: 	1142 
    -- CP-element group 603: successors 
    -- CP-element group 603:  members (5) 
      -- CP-element group 603: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_sample_completed_
      -- CP-element group 603: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Sample/$exit
      -- CP-element group 603: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Sample/word_access_start/$exit
      -- CP-element group 603: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Sample/word_access_start/word_0/$exit
      -- CP-element group 603: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Sample/word_access_start/word_0/ra
      -- 
    ra_8681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 603_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3852_load_0_ack_0, ack => zeropad3D_CP_2067_elements(603)); -- 
    -- CP-element group 604:  transition  input  output  bypass 
    -- CP-element group 604: predecessors 
    -- CP-element group 604: 	1142 
    -- CP-element group 604: successors 
    -- CP-element group 604: 	609 
    -- CP-element group 604:  members (12) 
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_update_completed_
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/$exit
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/word_access_complete/$exit
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/word_access_complete/word_0/$exit
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/word_access_complete/word_0/ca
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/LOAD_depth_high_3852_Merge/$entry
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/LOAD_depth_high_3852_Merge/$exit
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/LOAD_depth_high_3852_Merge/merge_req
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/LOAD_depth_high_3852_Merge/merge_ack
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_sample_start_
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_Sample/$entry
      -- CP-element group 604: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_Sample/rr
      -- 
    ca_8692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 604_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3852_load_0_ack_1, ack => zeropad3D_CP_2067_elements(604)); -- 
    rr_8771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(604), ack => type_cast_3862_inst_req_0); -- 
    -- CP-element group 605:  transition  input  bypass 
    -- CP-element group 605: predecessors 
    -- CP-element group 605: 	1142 
    -- CP-element group 605: successors 
    -- CP-element group 605:  members (5) 
      -- CP-element group 605: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_sample_completed_
      -- CP-element group 605: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Sample/$exit
      -- CP-element group 605: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Sample/word_access_start/$exit
      -- CP-element group 605: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Sample/word_access_start/word_0/$exit
      -- CP-element group 605: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Sample/word_access_start/word_0/ra
      -- 
    ra_8714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 605_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_3855_load_0_ack_0, ack => zeropad3D_CP_2067_elements(605)); -- 
    -- CP-element group 606:  fork  transition  input  output  bypass 
    -- CP-element group 606: predecessors 
    -- CP-element group 606: 	1142 
    -- CP-element group 606: successors 
    -- CP-element group 606: 	611 
    -- CP-element group 606: 	617 
    -- CP-element group 606:  members (15) 
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_Sample/rr
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_Sample/$entry
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_update_completed_
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/$exit
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/word_access_complete/$exit
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/word_access_complete/word_0/$exit
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/word_access_complete/word_0/ca
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/LOAD_out_depth_high_3855_Merge/$entry
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/LOAD_out_depth_high_3855_Merge/$exit
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/LOAD_out_depth_high_3855_Merge/merge_req
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/LOAD_out_depth_high_3855_Merge/merge_ack
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_sample_start_
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_Sample/$entry
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_Sample/rr
      -- CP-element group 606: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_sample_start_
      -- 
    ca_8725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 606_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_3855_load_0_ack_1, ack => zeropad3D_CP_2067_elements(606)); -- 
    rr_8785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(606), ack => type_cast_3866_inst_req_0); -- 
    rr_8827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(606), ack => type_cast_3883_inst_req_0); -- 
    -- CP-element group 607:  transition  input  bypass 
    -- CP-element group 607: predecessors 
    -- CP-element group 607: 	1142 
    -- CP-element group 607: successors 
    -- CP-element group 607:  members (5) 
      -- CP-element group 607: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_sample_completed_
      -- CP-element group 607: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Sample/$exit
      -- CP-element group 607: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Sample/word_access_start/$exit
      -- CP-element group 607: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Sample/word_access_start/word_0/$exit
      -- CP-element group 607: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Sample/word_access_start/word_0/ra
      -- 
    ra_8747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 607_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_3858_load_0_ack_0, ack => zeropad3D_CP_2067_elements(607)); -- 
    -- CP-element group 608:  transition  input  output  bypass 
    -- CP-element group 608: predecessors 
    -- CP-element group 608: 	1142 
    -- CP-element group 608: successors 
    -- CP-element group 608: 	613 
    -- CP-element group 608:  members (12) 
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_update_completed_
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/$exit
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/word_access_complete/$exit
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/word_access_complete/word_0/$exit
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/word_access_complete/word_0/ca
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/LOAD_out_col_high_3858_Merge/$entry
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/LOAD_out_col_high_3858_Merge/$exit
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/LOAD_out_col_high_3858_Merge/merge_req
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/LOAD_out_col_high_3858_Merge/merge_ack
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_sample_start_
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_Sample/$entry
      -- CP-element group 608: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_Sample/rr
      -- 
    ca_8758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 608_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_3858_load_0_ack_1, ack => zeropad3D_CP_2067_elements(608)); -- 
    rr_8799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(608), ack => type_cast_3870_inst_req_0); -- 
    -- CP-element group 609:  transition  input  bypass 
    -- CP-element group 609: predecessors 
    -- CP-element group 609: 	604 
    -- CP-element group 609: successors 
    -- CP-element group 609:  members (3) 
      -- CP-element group 609: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_sample_completed_
      -- CP-element group 609: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_Sample/$exit
      -- CP-element group 609: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_Sample/ra
      -- 
    ra_8772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 609_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3862_inst_ack_0, ack => zeropad3D_CP_2067_elements(609)); -- 
    -- CP-element group 610:  transition  input  bypass 
    -- CP-element group 610: predecessors 
    -- CP-element group 610: 	1142 
    -- CP-element group 610: successors 
    -- CP-element group 610: 	619 
    -- CP-element group 610:  members (3) 
      -- CP-element group 610: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_update_completed_
      -- CP-element group 610: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_Update/$exit
      -- CP-element group 610: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_Update/ca
      -- 
    ca_8777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 610_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3862_inst_ack_1, ack => zeropad3D_CP_2067_elements(610)); -- 
    -- CP-element group 611:  transition  input  bypass 
    -- CP-element group 611: predecessors 
    -- CP-element group 611: 	606 
    -- CP-element group 611: successors 
    -- CP-element group 611:  members (3) 
      -- CP-element group 611: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_sample_completed_
      -- CP-element group 611: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_Sample/$exit
      -- CP-element group 611: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_Sample/ra
      -- 
    ra_8786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 611_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3866_inst_ack_0, ack => zeropad3D_CP_2067_elements(611)); -- 
    -- CP-element group 612:  transition  input  bypass 
    -- CP-element group 612: predecessors 
    -- CP-element group 612: 	1142 
    -- CP-element group 612: successors 
    -- CP-element group 612: 	619 
    -- CP-element group 612:  members (3) 
      -- CP-element group 612: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_update_completed_
      -- CP-element group 612: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_Update/$exit
      -- CP-element group 612: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_Update/ca
      -- 
    ca_8791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 612_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3866_inst_ack_1, ack => zeropad3D_CP_2067_elements(612)); -- 
    -- CP-element group 613:  transition  input  bypass 
    -- CP-element group 613: predecessors 
    -- CP-element group 613: 	608 
    -- CP-element group 613: successors 
    -- CP-element group 613:  members (3) 
      -- CP-element group 613: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_sample_completed_
      -- CP-element group 613: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_Sample/$exit
      -- CP-element group 613: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_Sample/ra
      -- 
    ra_8800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 613_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3870_inst_ack_0, ack => zeropad3D_CP_2067_elements(613)); -- 
    -- CP-element group 614:  transition  input  bypass 
    -- CP-element group 614: predecessors 
    -- CP-element group 614: 	1142 
    -- CP-element group 614: successors 
    -- CP-element group 614: 	619 
    -- CP-element group 614:  members (3) 
      -- CP-element group 614: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_update_completed_
      -- CP-element group 614: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_Update/$exit
      -- CP-element group 614: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_Update/ca
      -- 
    ca_8805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 614_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3870_inst_ack_1, ack => zeropad3D_CP_2067_elements(614)); -- 
    -- CP-element group 615:  transition  input  bypass 
    -- CP-element group 615: predecessors 
    -- CP-element group 615: 	602 
    -- CP-element group 615: successors 
    -- CP-element group 615:  members (3) 
      -- CP-element group 615: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_sample_completed_
      -- CP-element group 615: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_Sample/$exit
      -- CP-element group 615: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_Sample/ra
      -- 
    ra_8814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 615_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3879_inst_ack_0, ack => zeropad3D_CP_2067_elements(615)); -- 
    -- CP-element group 616:  transition  input  bypass 
    -- CP-element group 616: predecessors 
    -- CP-element group 616: 	1142 
    -- CP-element group 616: successors 
    -- CP-element group 616: 	619 
    -- CP-element group 616:  members (3) 
      -- CP-element group 616: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_update_completed_
      -- CP-element group 616: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_Update/$exit
      -- CP-element group 616: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_Update/ca
      -- 
    ca_8819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 616_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3879_inst_ack_1, ack => zeropad3D_CP_2067_elements(616)); -- 
    -- CP-element group 617:  transition  input  bypass 
    -- CP-element group 617: predecessors 
    -- CP-element group 617: 	606 
    -- CP-element group 617: successors 
    -- CP-element group 617:  members (3) 
      -- CP-element group 617: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_Sample/ra
      -- CP-element group 617: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_Sample/$exit
      -- CP-element group 617: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_sample_completed_
      -- 
    ra_8828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 617_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3883_inst_ack_0, ack => zeropad3D_CP_2067_elements(617)); -- 
    -- CP-element group 618:  transition  input  bypass 
    -- CP-element group 618: predecessors 
    -- CP-element group 618: 	1142 
    -- CP-element group 618: successors 
    -- CP-element group 618: 	619 
    -- CP-element group 618:  members (3) 
      -- CP-element group 618: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_Update/ca
      -- CP-element group 618: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_Update/$exit
      -- CP-element group 618: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_update_completed_
      -- 
    ca_8833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 618_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3883_inst_ack_1, ack => zeropad3D_CP_2067_elements(618)); -- 
    -- CP-element group 619:  join  fork  transition  place  output  bypass 
    -- CP-element group 619: predecessors 
    -- CP-element group 619: 	600 
    -- CP-element group 619: 	610 
    -- CP-element group 619: 	612 
    -- CP-element group 619: 	614 
    -- CP-element group 619: 	616 
    -- CP-element group 619: 	618 
    -- CP-element group 619: successors 
    -- CP-element group 619: 	1153 
    -- CP-element group 619: 	1154 
    -- CP-element group 619: 	1155 
    -- CP-element group 619: 	1157 
    -- CP-element group 619:  members (16) 
      -- CP-element group 619: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925__exit__
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331
      -- CP-element group 619: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/$exit
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3928/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/Sample/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/Sample/rr
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/Update/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/Update/cr
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3941/$entry
      -- CP-element group 619: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/$entry
      -- 
    rr_13287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(619), ack => type_cast_3940_inst_req_0); -- 
    cr_13292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(619), ack => type_cast_3940_inst_req_1); -- 
    zeropad3D_cp_element_group_619: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_619"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(600) & zeropad3D_CP_2067_elements(610) & zeropad3D_CP_2067_elements(612) & zeropad3D_CP_2067_elements(614) & zeropad3D_CP_2067_elements(616) & zeropad3D_CP_2067_elements(618);
      gj_zeropad3D_cp_element_group_619 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(619), clk => clk, reset => reset); --
    end block;
    -- CP-element group 620:  transition  input  bypass 
    -- CP-element group 620: predecessors 
    -- CP-element group 620: 	1163 
    -- CP-element group 620: successors 
    -- CP-element group 620:  members (3) 
      -- CP-element group 620: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_Sample/ra
      -- CP-element group 620: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_Sample/$exit
      -- CP-element group 620: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_sample_completed_
      -- 
    ra_8845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 620_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3952_inst_ack_0, ack => zeropad3D_CP_2067_elements(620)); -- 
    -- CP-element group 621:  branch  transition  place  input  output  bypass 
    -- CP-element group 621: predecessors 
    -- CP-element group 621: 	1163 
    -- CP-element group 621: successors 
    -- CP-element group 621: 	622 
    -- CP-element group 621: 	623 
    -- CP-element group 621:  members (13) 
      -- CP-element group 621: 	 branch_block_stmt_655/if_stmt_3961__entry__
      -- CP-element group 621: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960__exit__
      -- CP-element group 621: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/$exit
      -- CP-element group 621: 	 branch_block_stmt_655/if_stmt_3961_else_link/$entry
      -- CP-element group 621: 	 branch_block_stmt_655/if_stmt_3961_if_link/$entry
      -- CP-element group 621: 	 branch_block_stmt_655/if_stmt_3961_eval_test/branch_req
      -- CP-element group 621: 	 branch_block_stmt_655/if_stmt_3961_eval_test/$exit
      -- CP-element group 621: 	 branch_block_stmt_655/if_stmt_3961_eval_test/$entry
      -- CP-element group 621: 	 branch_block_stmt_655/if_stmt_3961_dead_link/$entry
      -- CP-element group 621: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_Update/ca
      -- CP-element group 621: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_Update/$exit
      -- CP-element group 621: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_update_completed_
      -- CP-element group 621: 	 branch_block_stmt_655/R_cmp1336_3962_place
      -- 
    ca_8850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 621_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3952_inst_ack_1, ack => zeropad3D_CP_2067_elements(621)); -- 
    branch_req_8858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(621), ack => if_stmt_3961_branch_req_0); -- 
    -- CP-element group 622:  transition  place  input  bypass 
    -- CP-element group 622: predecessors 
    -- CP-element group 622: 	621 
    -- CP-element group 622: successors 
    -- CP-element group 622: 	1164 
    -- CP-element group 622:  members (5) 
      -- CP-element group 622: 	 branch_block_stmt_655/if_stmt_3961_if_link/if_choice_transition
      -- CP-element group 622: 	 branch_block_stmt_655/if_stmt_3961_if_link/$exit
      -- CP-element group 622: 	 branch_block_stmt_655/whilex_xbody1331_ifx_xthen1366
      -- CP-element group 622: 	 branch_block_stmt_655/whilex_xbody1331_ifx_xthen1366_PhiReq/$entry
      -- CP-element group 622: 	 branch_block_stmt_655/whilex_xbody1331_ifx_xthen1366_PhiReq/$exit
      -- 
    if_choice_transition_8863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 622_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3961_branch_ack_1, ack => zeropad3D_CP_2067_elements(622)); -- 
    -- CP-element group 623:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 623: predecessors 
    -- CP-element group 623: 	621 
    -- CP-element group 623: successors 
    -- CP-element group 623: 	624 
    -- CP-element group 623: 	625 
    -- CP-element group 623: 	627 
    -- CP-element group 623:  members (27) 
      -- CP-element group 623: 	 branch_block_stmt_655/merge_stmt_3967__exit__
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986__entry__
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Sample/word_access_start/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Sample/word_access_start/word_0/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Sample/word_access_start/word_0/rr
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Sample/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_Update/cr
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_Update/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/if_stmt_3961_else_link/else_choice_transition
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_root_address_calculated
      -- CP-element group 623: 	 branch_block_stmt_655/if_stmt_3961_else_link/$exit
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_word_address_calculated
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_update_start_
      -- CP-element group 623: 	 branch_block_stmt_655/whilex_xbody1331_lorx_xlhsx_xfalse1338
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_update_start_
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/word_access_complete/word_0/cr
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/word_access_complete/word_0/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_sample_start_
      -- CP-element group 623: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/word_access_complete/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/whilex_xbody1331_lorx_xlhsx_xfalse1338_PhiReq/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/whilex_xbody1331_lorx_xlhsx_xfalse1338_PhiReq/$exit
      -- CP-element group 623: 	 branch_block_stmt_655/merge_stmt_3967_PhiReqMerge
      -- CP-element group 623: 	 branch_block_stmt_655/merge_stmt_3967_PhiAck/$entry
      -- CP-element group 623: 	 branch_block_stmt_655/merge_stmt_3967_PhiAck/$exit
      -- CP-element group 623: 	 branch_block_stmt_655/merge_stmt_3967_PhiAck/dummy
      -- 
    else_choice_transition_8867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 623_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3961_branch_ack_0, ack => zeropad3D_CP_2067_elements(623)); -- 
    rr_8888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(623), ack => LOAD_row_high_3969_load_0_req_0); -- 
    cr_8918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(623), ack => type_cast_3973_inst_req_1); -- 
    cr_8899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(623), ack => LOAD_row_high_3969_load_0_req_1); -- 
    -- CP-element group 624:  transition  input  bypass 
    -- CP-element group 624: predecessors 
    -- CP-element group 624: 	623 
    -- CP-element group 624: successors 
    -- CP-element group 624:  members (5) 
      -- CP-element group 624: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Sample/$exit
      -- CP-element group 624: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Sample/word_access_start/$exit
      -- CP-element group 624: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Sample/word_access_start/word_0/$exit
      -- CP-element group 624: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Sample/word_access_start/word_0/ra
      -- CP-element group 624: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_sample_completed_
      -- 
    ra_8889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 624_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3969_load_0_ack_0, ack => zeropad3D_CP_2067_elements(624)); -- 
    -- CP-element group 625:  transition  input  output  bypass 
    -- CP-element group 625: predecessors 
    -- CP-element group 625: 	623 
    -- CP-element group 625: successors 
    -- CP-element group 625: 	626 
    -- CP-element group 625:  members (12) 
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_Sample/rr
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_Sample/$entry
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_update_completed_
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_sample_start_
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/LOAD_row_high_3969_Merge/merge_ack
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/LOAD_row_high_3969_Merge/merge_req
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/LOAD_row_high_3969_Merge/$exit
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/LOAD_row_high_3969_Merge/$entry
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/word_access_complete/word_0/ca
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/word_access_complete/word_0/$exit
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/word_access_complete/$exit
      -- CP-element group 625: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/LOAD_row_high_3969_Update/$exit
      -- 
    ca_8900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 625_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3969_load_0_ack_1, ack => zeropad3D_CP_2067_elements(625)); -- 
    rr_8913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(625), ack => type_cast_3973_inst_req_0); -- 
    -- CP-element group 626:  transition  input  bypass 
    -- CP-element group 626: predecessors 
    -- CP-element group 626: 	625 
    -- CP-element group 626: successors 
    -- CP-element group 626:  members (3) 
      -- CP-element group 626: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_Sample/ra
      -- CP-element group 626: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_Sample/$exit
      -- CP-element group 626: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_sample_completed_
      -- 
    ra_8914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 626_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3973_inst_ack_0, ack => zeropad3D_CP_2067_elements(626)); -- 
    -- CP-element group 627:  branch  transition  place  input  output  bypass 
    -- CP-element group 627: predecessors 
    -- CP-element group 627: 	623 
    -- CP-element group 627: successors 
    -- CP-element group 627: 	628 
    -- CP-element group 627: 	629 
    -- CP-element group 627:  members (13) 
      -- CP-element group 627: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986__exit__
      -- CP-element group 627: 	 branch_block_stmt_655/if_stmt_3987__entry__
      -- CP-element group 627: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_Update/ca
      -- CP-element group 627: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/$exit
      -- CP-element group 627: 	 branch_block_stmt_655/if_stmt_3987_dead_link/$entry
      -- CP-element group 627: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_Update/$exit
      -- CP-element group 627: 	 branch_block_stmt_655/R_cmp1346_3988_place
      -- CP-element group 627: 	 branch_block_stmt_655/assign_stmt_3970_to_assign_stmt_3986/type_cast_3973_update_completed_
      -- CP-element group 627: 	 branch_block_stmt_655/if_stmt_3987_else_link/$entry
      -- CP-element group 627: 	 branch_block_stmt_655/if_stmt_3987_if_link/$entry
      -- CP-element group 627: 	 branch_block_stmt_655/if_stmt_3987_eval_test/branch_req
      -- CP-element group 627: 	 branch_block_stmt_655/if_stmt_3987_eval_test/$exit
      -- CP-element group 627: 	 branch_block_stmt_655/if_stmt_3987_eval_test/$entry
      -- 
    ca_8919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 627_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3973_inst_ack_1, ack => zeropad3D_CP_2067_elements(627)); -- 
    branch_req_8927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(627), ack => if_stmt_3987_branch_req_0); -- 
    -- CP-element group 628:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 628: predecessors 
    -- CP-element group 628: 	627 
    -- CP-element group 628: successors 
    -- CP-element group 628: 	630 
    -- CP-element group 628: 	631 
    -- CP-element group 628:  members (18) 
      -- CP-element group 628: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005__entry__
      -- CP-element group 628: 	 branch_block_stmt_655/merge_stmt_3993__exit__
      -- CP-element group 628: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1338_lorx_xlhsx_xfalse1348
      -- CP-element group 628: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_Update/cr
      -- CP-element group 628: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_Update/$entry
      -- CP-element group 628: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_Sample/rr
      -- CP-element group 628: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_Sample/$entry
      -- CP-element group 628: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_update_start_
      -- CP-element group 628: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_sample_start_
      -- CP-element group 628: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/$entry
      -- CP-element group 628: 	 branch_block_stmt_655/if_stmt_3987_if_link/if_choice_transition
      -- CP-element group 628: 	 branch_block_stmt_655/if_stmt_3987_if_link/$exit
      -- CP-element group 628: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1338_lorx_xlhsx_xfalse1348_PhiReq/$entry
      -- CP-element group 628: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1338_lorx_xlhsx_xfalse1348_PhiReq/$exit
      -- CP-element group 628: 	 branch_block_stmt_655/merge_stmt_3993_PhiReqMerge
      -- CP-element group 628: 	 branch_block_stmt_655/merge_stmt_3993_PhiAck/$entry
      -- CP-element group 628: 	 branch_block_stmt_655/merge_stmt_3993_PhiAck/$exit
      -- CP-element group 628: 	 branch_block_stmt_655/merge_stmt_3993_PhiAck/dummy
      -- 
    if_choice_transition_8932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 628_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3987_branch_ack_1, ack => zeropad3D_CP_2067_elements(628)); -- 
    cr_8954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(628), ack => type_cast_3997_inst_req_1); -- 
    rr_8949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(628), ack => type_cast_3997_inst_req_0); -- 
    -- CP-element group 629:  transition  place  input  bypass 
    -- CP-element group 629: predecessors 
    -- CP-element group 629: 	627 
    -- CP-element group 629: successors 
    -- CP-element group 629: 	1164 
    -- CP-element group 629:  members (5) 
      -- CP-element group 629: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1338_ifx_xthen1366
      -- CP-element group 629: 	 branch_block_stmt_655/if_stmt_3987_else_link/else_choice_transition
      -- CP-element group 629: 	 branch_block_stmt_655/if_stmt_3987_else_link/$exit
      -- CP-element group 629: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1338_ifx_xthen1366_PhiReq/$entry
      -- CP-element group 629: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1338_ifx_xthen1366_PhiReq/$exit
      -- 
    else_choice_transition_8936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 629_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3987_branch_ack_0, ack => zeropad3D_CP_2067_elements(629)); -- 
    -- CP-element group 630:  transition  input  bypass 
    -- CP-element group 630: predecessors 
    -- CP-element group 630: 	628 
    -- CP-element group 630: successors 
    -- CP-element group 630:  members (3) 
      -- CP-element group 630: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_Sample/ra
      -- CP-element group 630: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_Sample/$exit
      -- CP-element group 630: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_sample_completed_
      -- 
    ra_8950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 630_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3997_inst_ack_0, ack => zeropad3D_CP_2067_elements(630)); -- 
    -- CP-element group 631:  branch  transition  place  input  output  bypass 
    -- CP-element group 631: predecessors 
    -- CP-element group 631: 	628 
    -- CP-element group 631: successors 
    -- CP-element group 631: 	632 
    -- CP-element group 631: 	633 
    -- CP-element group 631:  members (13) 
      -- CP-element group 631: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005__exit__
      -- CP-element group 631: 	 branch_block_stmt_655/if_stmt_4006__entry__
      -- CP-element group 631: 	 branch_block_stmt_655/if_stmt_4006_else_link/$entry
      -- CP-element group 631: 	 branch_block_stmt_655/if_stmt_4006_if_link/$entry
      -- CP-element group 631: 	 branch_block_stmt_655/R_cmp1353_4007_place
      -- CP-element group 631: 	 branch_block_stmt_655/if_stmt_4006_eval_test/branch_req
      -- CP-element group 631: 	 branch_block_stmt_655/if_stmt_4006_eval_test/$exit
      -- CP-element group 631: 	 branch_block_stmt_655/if_stmt_4006_eval_test/$entry
      -- CP-element group 631: 	 branch_block_stmt_655/if_stmt_4006_dead_link/$entry
      -- CP-element group 631: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_Update/ca
      -- CP-element group 631: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_Update/$exit
      -- CP-element group 631: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/type_cast_3997_update_completed_
      -- CP-element group 631: 	 branch_block_stmt_655/assign_stmt_3998_to_assign_stmt_4005/$exit
      -- 
    ca_8955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 631_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3997_inst_ack_1, ack => zeropad3D_CP_2067_elements(631)); -- 
    branch_req_8963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(631), ack => if_stmt_4006_branch_req_0); -- 
    -- CP-element group 632:  transition  place  input  bypass 
    -- CP-element group 632: predecessors 
    -- CP-element group 632: 	631 
    -- CP-element group 632: successors 
    -- CP-element group 632: 	1164 
    -- CP-element group 632:  members (5) 
      -- CP-element group 632: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1348_ifx_xthen1366
      -- CP-element group 632: 	 branch_block_stmt_655/if_stmt_4006_if_link/if_choice_transition
      -- CP-element group 632: 	 branch_block_stmt_655/if_stmt_4006_if_link/$exit
      -- CP-element group 632: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1348_ifx_xthen1366_PhiReq/$entry
      -- CP-element group 632: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1348_ifx_xthen1366_PhiReq/$exit
      -- 
    if_choice_transition_8968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 632_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4006_branch_ack_1, ack => zeropad3D_CP_2067_elements(632)); -- 
    -- CP-element group 633:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 633: predecessors 
    -- CP-element group 633: 	631 
    -- CP-element group 633: successors 
    -- CP-element group 633: 	634 
    -- CP-element group 633: 	635 
    -- CP-element group 633: 	637 
    -- CP-element group 633:  members (27) 
      -- CP-element group 633: 	 branch_block_stmt_655/merge_stmt_4012__exit__
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037__entry__
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_update_start_
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_Update/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_Update/cr
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/word_access_complete/word_0/cr
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/word_access_complete/word_0/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/word_access_complete/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Sample/word_access_start/word_0/rr
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Sample/word_access_start/word_0/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Sample/word_access_start/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Sample/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_root_address_calculated
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_word_address_calculated
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_update_start_
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_sample_start_
      -- CP-element group 633: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1355
      -- CP-element group 633: 	 branch_block_stmt_655/if_stmt_4006_else_link/else_choice_transition
      -- CP-element group 633: 	 branch_block_stmt_655/if_stmt_4006_else_link/$exit
      -- CP-element group 633: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1355_PhiReq/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1355_PhiReq/$exit
      -- CP-element group 633: 	 branch_block_stmt_655/merge_stmt_4012_PhiReqMerge
      -- CP-element group 633: 	 branch_block_stmt_655/merge_stmt_4012_PhiAck/$entry
      -- CP-element group 633: 	 branch_block_stmt_655/merge_stmt_4012_PhiAck/$exit
      -- CP-element group 633: 	 branch_block_stmt_655/merge_stmt_4012_PhiAck/dummy
      -- 
    else_choice_transition_8972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 633_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4006_branch_ack_0, ack => zeropad3D_CP_2067_elements(633)); -- 
    cr_9023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(633), ack => type_cast_4018_inst_req_1); -- 
    cr_9004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(633), ack => LOAD_col_high_4014_load_0_req_1); -- 
    rr_8993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(633), ack => LOAD_col_high_4014_load_0_req_0); -- 
    -- CP-element group 634:  transition  input  bypass 
    -- CP-element group 634: predecessors 
    -- CP-element group 634: 	633 
    -- CP-element group 634: successors 
    -- CP-element group 634:  members (5) 
      -- CP-element group 634: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Sample/word_access_start/word_0/ra
      -- CP-element group 634: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Sample/word_access_start/word_0/$exit
      -- CP-element group 634: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Sample/word_access_start/$exit
      -- CP-element group 634: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Sample/$exit
      -- CP-element group 634: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_sample_completed_
      -- 
    ra_8994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 634_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4014_load_0_ack_0, ack => zeropad3D_CP_2067_elements(634)); -- 
    -- CP-element group 635:  transition  input  output  bypass 
    -- CP-element group 635: predecessors 
    -- CP-element group 635: 	633 
    -- CP-element group 635: successors 
    -- CP-element group 635: 	636 
    -- CP-element group 635:  members (12) 
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_Sample/$entry
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_Sample/rr
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_sample_start_
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/LOAD_col_high_4014_Merge/merge_ack
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/LOAD_col_high_4014_Merge/merge_req
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/LOAD_col_high_4014_Merge/$exit
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/LOAD_col_high_4014_Merge/$entry
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/word_access_complete/word_0/ca
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/word_access_complete/word_0/$exit
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/word_access_complete/$exit
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_Update/$exit
      -- CP-element group 635: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/LOAD_col_high_4014_update_completed_
      -- 
    ca_9005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 635_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4014_load_0_ack_1, ack => zeropad3D_CP_2067_elements(635)); -- 
    rr_9018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(635), ack => type_cast_4018_inst_req_0); -- 
    -- CP-element group 636:  transition  input  bypass 
    -- CP-element group 636: predecessors 
    -- CP-element group 636: 	635 
    -- CP-element group 636: successors 
    -- CP-element group 636:  members (3) 
      -- CP-element group 636: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_sample_completed_
      -- CP-element group 636: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_Sample/$exit
      -- CP-element group 636: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_Sample/ra
      -- 
    ra_9019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 636_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4018_inst_ack_0, ack => zeropad3D_CP_2067_elements(636)); -- 
    -- CP-element group 637:  branch  transition  place  input  output  bypass 
    -- CP-element group 637: predecessors 
    -- CP-element group 637: 	633 
    -- CP-element group 637: successors 
    -- CP-element group 637: 	638 
    -- CP-element group 637: 	639 
    -- CP-element group 637:  members (13) 
      -- CP-element group 637: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037__exit__
      -- CP-element group 637: 	 branch_block_stmt_655/if_stmt_4038__entry__
      -- CP-element group 637: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_update_completed_
      -- CP-element group 637: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_Update/$exit
      -- CP-element group 637: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/type_cast_4018_Update/ca
      -- CP-element group 637: 	 branch_block_stmt_655/if_stmt_4038_else_link/$entry
      -- CP-element group 637: 	 branch_block_stmt_655/assign_stmt_4015_to_assign_stmt_4037/$exit
      -- CP-element group 637: 	 branch_block_stmt_655/if_stmt_4038_if_link/$entry
      -- CP-element group 637: 	 branch_block_stmt_655/R_cmp1364_4039_place
      -- CP-element group 637: 	 branch_block_stmt_655/if_stmt_4038_eval_test/branch_req
      -- CP-element group 637: 	 branch_block_stmt_655/if_stmt_4038_eval_test/$exit
      -- CP-element group 637: 	 branch_block_stmt_655/if_stmt_4038_eval_test/$entry
      -- CP-element group 637: 	 branch_block_stmt_655/if_stmt_4038_dead_link/$entry
      -- 
    ca_9024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 637_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4018_inst_ack_1, ack => zeropad3D_CP_2067_elements(637)); -- 
    branch_req_9032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(637), ack => if_stmt_4038_branch_req_0); -- 
    -- CP-element group 638:  fork  transition  place  input  output  bypass 
    -- CP-element group 638: predecessors 
    -- CP-element group 638: 	637 
    -- CP-element group 638: successors 
    -- CP-element group 638: 	654 
    -- CP-element group 638: 	655 
    -- CP-element group 638: 	657 
    -- CP-element group 638: 	659 
    -- CP-element group 638: 	661 
    -- CP-element group 638: 	663 
    -- CP-element group 638: 	665 
    -- CP-element group 638: 	667 
    -- CP-element group 638: 	669 
    -- CP-element group 638: 	672 
    -- CP-element group 638:  members (46) 
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207__entry__
      -- CP-element group 638: 	 branch_block_stmt_655/merge_stmt_4102__exit__
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_complete/req
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_Update/req
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_Sample/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_Update/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_update_start_
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_sample_start_
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_Update/cr
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_update_start_
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_update_start
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_Update/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1355_ifx_xelse1387
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_complete/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/if_stmt_4038_if_link/if_choice_transition
      -- CP-element group 638: 	 branch_block_stmt_655/if_stmt_4038_if_link/$exit
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_update_start_
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_Update/cr
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_Update/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_update_start_
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_Sample/rr
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/word_access_complete/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/word_access_complete/word_0/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/word_access_complete/word_0/cr
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_update_start_
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_Update/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_Update/cr
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_update_start_
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_update_start
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_Update/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_Update/req
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_complete/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_complete/req
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_update_start_
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Update/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Update/word_access_complete/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Update/word_access_complete/word_0/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Update/word_access_complete/word_0/cr
      -- CP-element group 638: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1355_ifx_xelse1387_PhiReq/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1355_ifx_xelse1387_PhiReq/$exit
      -- CP-element group 638: 	 branch_block_stmt_655/merge_stmt_4102_PhiReqMerge
      -- CP-element group 638: 	 branch_block_stmt_655/merge_stmt_4102_PhiAck/$entry
      -- CP-element group 638: 	 branch_block_stmt_655/merge_stmt_4102_PhiAck/$exit
      -- CP-element group 638: 	 branch_block_stmt_655/merge_stmt_4102_PhiAck/dummy
      -- 
    if_choice_transition_9037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 638_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4038_branch_ack_1, ack => zeropad3D_CP_2067_elements(638)); -- 
    req_9260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => addr_of_4177_final_reg_req_1); -- 
    req_9245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => array_obj_ref_4176_index_offset_req_1); -- 
    cr_9214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => type_cast_4170_inst_req_1); -- 
    cr_9200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => type_cast_4106_inst_req_1); -- 
    rr_9195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => type_cast_4106_inst_req_0); -- 
    cr_9305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => ptr_deref_4181_load_0_req_1); -- 
    cr_9324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => type_cast_4195_inst_req_1); -- 
    req_9355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => array_obj_ref_4201_index_offset_req_1); -- 
    req_9370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => addr_of_4202_final_reg_req_1); -- 
    cr_9420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(638), ack => ptr_deref_4205_store_0_req_1); -- 
    -- CP-element group 639:  transition  place  input  bypass 
    -- CP-element group 639: predecessors 
    -- CP-element group 639: 	637 
    -- CP-element group 639: successors 
    -- CP-element group 639: 	1164 
    -- CP-element group 639:  members (5) 
      -- CP-element group 639: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1355_ifx_xthen1366
      -- CP-element group 639: 	 branch_block_stmt_655/if_stmt_4038_else_link/else_choice_transition
      -- CP-element group 639: 	 branch_block_stmt_655/if_stmt_4038_else_link/$exit
      -- CP-element group 639: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1355_ifx_xthen1366_PhiReq/$entry
      -- CP-element group 639: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1355_ifx_xthen1366_PhiReq/$exit
      -- 
    else_choice_transition_9041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 639_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4038_branch_ack_0, ack => zeropad3D_CP_2067_elements(639)); -- 
    -- CP-element group 640:  transition  input  bypass 
    -- CP-element group 640: predecessors 
    -- CP-element group 640: 	1164 
    -- CP-element group 640: successors 
    -- CP-element group 640:  members (3) 
      -- CP-element group 640: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_Sample/ra
      -- CP-element group 640: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_Sample/$exit
      -- CP-element group 640: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_sample_completed_
      -- 
    ra_9055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 640_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4048_inst_ack_0, ack => zeropad3D_CP_2067_elements(640)); -- 
    -- CP-element group 641:  transition  input  bypass 
    -- CP-element group 641: predecessors 
    -- CP-element group 641: 	1164 
    -- CP-element group 641: successors 
    -- CP-element group 641: 	644 
    -- CP-element group 641:  members (3) 
      -- CP-element group 641: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_Update/$exit
      -- CP-element group 641: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_update_completed_
      -- CP-element group 641: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_Update/ca
      -- 
    ca_9060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 641_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4048_inst_ack_1, ack => zeropad3D_CP_2067_elements(641)); -- 
    -- CP-element group 642:  transition  input  bypass 
    -- CP-element group 642: predecessors 
    -- CP-element group 642: 	1164 
    -- CP-element group 642: successors 
    -- CP-element group 642:  members (3) 
      -- CP-element group 642: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_Sample/ra
      -- CP-element group 642: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_Sample/$exit
      -- CP-element group 642: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_sample_completed_
      -- 
    ra_9069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 642_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4053_inst_ack_0, ack => zeropad3D_CP_2067_elements(642)); -- 
    -- CP-element group 643:  transition  input  bypass 
    -- CP-element group 643: predecessors 
    -- CP-element group 643: 	1164 
    -- CP-element group 643: successors 
    -- CP-element group 643: 	644 
    -- CP-element group 643:  members (3) 
      -- CP-element group 643: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_Update/ca
      -- CP-element group 643: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_Update/$exit
      -- CP-element group 643: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_update_completed_
      -- 
    ca_9074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 643_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4053_inst_ack_1, ack => zeropad3D_CP_2067_elements(643)); -- 
    -- CP-element group 644:  join  transition  output  bypass 
    -- CP-element group 644: predecessors 
    -- CP-element group 644: 	641 
    -- CP-element group 644: 	643 
    -- CP-element group 644: successors 
    -- CP-element group 644: 	645 
    -- CP-element group 644:  members (3) 
      -- CP-element group 644: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_Sample/rr
      -- CP-element group 644: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_Sample/$entry
      -- CP-element group 644: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_sample_start_
      -- 
    rr_9082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(644), ack => type_cast_4087_inst_req_0); -- 
    zeropad3D_cp_element_group_644: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_644"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(641) & zeropad3D_CP_2067_elements(643);
      gj_zeropad3D_cp_element_group_644 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(644), clk => clk, reset => reset); --
    end block;
    -- CP-element group 645:  transition  input  bypass 
    -- CP-element group 645: predecessors 
    -- CP-element group 645: 	644 
    -- CP-element group 645: successors 
    -- CP-element group 645:  members (3) 
      -- CP-element group 645: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_Sample/ra
      -- CP-element group 645: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_Sample/$exit
      -- CP-element group 645: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_sample_completed_
      -- 
    ra_9083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 645_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4087_inst_ack_0, ack => zeropad3D_CP_2067_elements(645)); -- 
    -- CP-element group 646:  transition  input  output  bypass 
    -- CP-element group 646: predecessors 
    -- CP-element group 646: 	1164 
    -- CP-element group 646: successors 
    -- CP-element group 646: 	647 
    -- CP-element group 646:  members (16) 
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_resized_1
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_scaled_1
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_Update/ca
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_Update/$exit
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_update_completed_
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_Sample/req
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_Sample/$entry
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_scale_1/scale_rename_ack
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_scale_1/scale_rename_req
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_scale_1/$exit
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_scale_1/$entry
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_resize_1/index_resize_ack
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_resize_1/index_resize_req
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_resize_1/$exit
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_resize_1/$entry
      -- CP-element group 646: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_index_computed_1
      -- 
    ca_9088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 646_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4087_inst_ack_1, ack => zeropad3D_CP_2067_elements(646)); -- 
    req_9113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(646), ack => array_obj_ref_4093_index_offset_req_0); -- 
    -- CP-element group 647:  transition  input  bypass 
    -- CP-element group 647: predecessors 
    -- CP-element group 647: 	646 
    -- CP-element group 647: successors 
    -- CP-element group 647: 	653 
    -- CP-element group 647:  members (3) 
      -- CP-element group 647: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_Sample/ack
      -- CP-element group 647: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_Sample/$exit
      -- CP-element group 647: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_sample_complete
      -- 
    ack_9114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 647_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4093_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(647)); -- 
    -- CP-element group 648:  transition  input  output  bypass 
    -- CP-element group 648: predecessors 
    -- CP-element group 648: 	1164 
    -- CP-element group 648: successors 
    -- CP-element group 648: 	649 
    -- CP-element group 648:  members (11) 
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_offset_calculated
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_root_address_calculated
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_request/req
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_request/$entry
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_sample_start_
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_base_plus_offset/sum_rename_ack
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_base_plus_offset/sum_rename_req
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_base_plus_offset/$exit
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_base_plus_offset/$entry
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_Update/ack
      -- CP-element group 648: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_Update/$exit
      -- 
    ack_9119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 648_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4093_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(648)); -- 
    req_9128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(648), ack => addr_of_4094_final_reg_req_0); -- 
    -- CP-element group 649:  transition  input  bypass 
    -- CP-element group 649: predecessors 
    -- CP-element group 649: 	648 
    -- CP-element group 649: successors 
    -- CP-element group 649:  members (3) 
      -- CP-element group 649: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_request/ack
      -- CP-element group 649: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_request/$exit
      -- CP-element group 649: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_sample_completed_
      -- 
    ack_9129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 649_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4094_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(649)); -- 
    -- CP-element group 650:  join  fork  transition  input  output  bypass 
    -- CP-element group 650: predecessors 
    -- CP-element group 650: 	1164 
    -- CP-element group 650: successors 
    -- CP-element group 650: 	651 
    -- CP-element group 650:  members (28) 
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_root_address_calculated
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_sample_start_
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_addr_resize/$exit
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_addr_resize/base_resize_ack
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_complete/ack
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_update_completed_
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_complete/$exit
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_addr_resize/base_resize_req
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_word_address_calculated
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_addr_resize/$entry
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_address_resized
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/word_access_start/word_0/rr
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/word_access_start/word_0/$entry
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/word_access_start/$entry
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/ptr_deref_4097_Split/split_ack
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/ptr_deref_4097_Split/split_req
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/ptr_deref_4097_Split/$exit
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/ptr_deref_4097_Split/$entry
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/$entry
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_word_addrgen/root_register_ack
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_word_addrgen/root_register_req
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_address_calculated
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_word_addrgen/$exit
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_word_addrgen/$entry
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_plus_offset/sum_rename_ack
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_plus_offset/sum_rename_req
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_plus_offset/$exit
      -- CP-element group 650: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_base_plus_offset/$entry
      -- 
    ack_9134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 650_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4094_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(650)); -- 
    rr_9172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(650), ack => ptr_deref_4097_store_0_req_0); -- 
    -- CP-element group 651:  transition  input  bypass 
    -- CP-element group 651: predecessors 
    -- CP-element group 651: 	650 
    -- CP-element group 651: successors 
    -- CP-element group 651:  members (5) 
      -- CP-element group 651: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/word_access_start/word_0/ra
      -- CP-element group 651: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/word_access_start/word_0/$exit
      -- CP-element group 651: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/word_access_start/$exit
      -- CP-element group 651: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Sample/$exit
      -- CP-element group 651: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_sample_completed_
      -- 
    ra_9173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 651_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4097_store_0_ack_0, ack => zeropad3D_CP_2067_elements(651)); -- 
    -- CP-element group 652:  transition  input  bypass 
    -- CP-element group 652: predecessors 
    -- CP-element group 652: 	1164 
    -- CP-element group 652: successors 
    -- CP-element group 652: 	653 
    -- CP-element group 652:  members (5) 
      -- CP-element group 652: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Update/word_access_complete/word_0/ca
      -- CP-element group 652: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Update/word_access_complete/word_0/$exit
      -- CP-element group 652: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Update/word_access_complete/$exit
      -- CP-element group 652: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Update/$exit
      -- CP-element group 652: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_update_completed_
      -- 
    ca_9184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 652_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4097_store_0_ack_1, ack => zeropad3D_CP_2067_elements(652)); -- 
    -- CP-element group 653:  join  transition  place  bypass 
    -- CP-element group 653: predecessors 
    -- CP-element group 653: 	647 
    -- CP-element group 653: 	652 
    -- CP-element group 653: successors 
    -- CP-element group 653: 	1165 
    -- CP-element group 653:  members (5) 
      -- CP-element group 653: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100__exit__
      -- CP-element group 653: 	 branch_block_stmt_655/ifx_xthen1366_ifx_xend1435
      -- CP-element group 653: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/$exit
      -- CP-element group 653: 	 branch_block_stmt_655/ifx_xthen1366_ifx_xend1435_PhiReq/$entry
      -- CP-element group 653: 	 branch_block_stmt_655/ifx_xthen1366_ifx_xend1435_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_653: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_653"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(647) & zeropad3D_CP_2067_elements(652);
      gj_zeropad3D_cp_element_group_653 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(653), clk => clk, reset => reset); --
    end block;
    -- CP-element group 654:  transition  input  bypass 
    -- CP-element group 654: predecessors 
    -- CP-element group 654: 	638 
    -- CP-element group 654: successors 
    -- CP-element group 654:  members (3) 
      -- CP-element group 654: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_Sample/$exit
      -- CP-element group 654: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_sample_completed_
      -- CP-element group 654: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_Sample/ra
      -- 
    ra_9196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 654_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4106_inst_ack_0, ack => zeropad3D_CP_2067_elements(654)); -- 
    -- CP-element group 655:  fork  transition  input  output  bypass 
    -- CP-element group 655: predecessors 
    -- CP-element group 655: 	638 
    -- CP-element group 655: successors 
    -- CP-element group 655: 	656 
    -- CP-element group 655: 	664 
    -- CP-element group 655:  members (9) 
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_update_completed_
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_Sample/rr
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_Sample/$entry
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_sample_start_
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_Update/ca
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4106_Update/$exit
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_sample_start_
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_Sample/$entry
      -- CP-element group 655: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_Sample/rr
      -- 
    ca_9201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 655_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4106_inst_ack_1, ack => zeropad3D_CP_2067_elements(655)); -- 
    rr_9209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(655), ack => type_cast_4170_inst_req_0); -- 
    rr_9319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(655), ack => type_cast_4195_inst_req_0); -- 
    -- CP-element group 656:  transition  input  bypass 
    -- CP-element group 656: predecessors 
    -- CP-element group 656: 	655 
    -- CP-element group 656: successors 
    -- CP-element group 656:  members (3) 
      -- CP-element group 656: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_Sample/ra
      -- CP-element group 656: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_Sample/$exit
      -- CP-element group 656: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_sample_completed_
      -- 
    ra_9210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 656_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4170_inst_ack_0, ack => zeropad3D_CP_2067_elements(656)); -- 
    -- CP-element group 657:  transition  input  output  bypass 
    -- CP-element group 657: predecessors 
    -- CP-element group 657: 	638 
    -- CP-element group 657: successors 
    -- CP-element group 657: 	658 
    -- CP-element group 657:  members (16) 
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_Update/ca
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_Sample/req
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_Update/$exit
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_Sample/$entry
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_scale_1/scale_rename_ack
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_scale_1/scale_rename_req
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_scale_1/$exit
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_scale_1/$entry
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_resize_1/index_resize_ack
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_resize_1/index_resize_req
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_resize_1/$exit
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_resize_1/$entry
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4170_update_completed_
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_computed_1
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_scaled_1
      -- CP-element group 657: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_index_resized_1
      -- 
    ca_9215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 657_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4170_inst_ack_1, ack => zeropad3D_CP_2067_elements(657)); -- 
    req_9240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(657), ack => array_obj_ref_4176_index_offset_req_0); -- 
    -- CP-element group 658:  transition  input  bypass 
    -- CP-element group 658: predecessors 
    -- CP-element group 658: 	657 
    -- CP-element group 658: successors 
    -- CP-element group 658: 	673 
    -- CP-element group 658:  members (3) 
      -- CP-element group 658: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_Sample/ack
      -- CP-element group 658: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_Sample/$exit
      -- CP-element group 658: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_sample_complete
      -- 
    ack_9241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 658_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4176_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(658)); -- 
    -- CP-element group 659:  transition  input  output  bypass 
    -- CP-element group 659: predecessors 
    -- CP-element group 659: 	638 
    -- CP-element group 659: successors 
    -- CP-element group 659: 	660 
    -- CP-element group 659:  members (11) 
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_request/$entry
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_sample_start_
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_Update/$exit
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_base_plus_offset/sum_rename_ack
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_base_plus_offset/sum_rename_req
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_base_plus_offset/$exit
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_base_plus_offset/$entry
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_request/req
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_final_index_sum_regn_Update/ack
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_offset_calculated
      -- CP-element group 659: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4176_root_address_calculated
      -- 
    ack_9246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 659_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4176_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(659)); -- 
    req_9255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(659), ack => addr_of_4177_final_reg_req_0); -- 
    -- CP-element group 660:  transition  input  bypass 
    -- CP-element group 660: predecessors 
    -- CP-element group 660: 	659 
    -- CP-element group 660: successors 
    -- CP-element group 660:  members (3) 
      -- CP-element group 660: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_sample_completed_
      -- CP-element group 660: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_request/ack
      -- CP-element group 660: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_request/$exit
      -- 
    ack_9256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 660_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4177_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(660)); -- 
    -- CP-element group 661:  join  fork  transition  input  output  bypass 
    -- CP-element group 661: predecessors 
    -- CP-element group 661: 	638 
    -- CP-element group 661: successors 
    -- CP-element group 661: 	662 
    -- CP-element group 661:  members (24) 
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_address_calculated
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_complete/$exit
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_root_address_calculated
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_sample_start_
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_address_resized
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_word_address_calculated
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_complete/ack
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4177_update_completed_
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_addr_resize/$entry
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_addr_resize/$exit
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_addr_resize/base_resize_req
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_addr_resize/base_resize_ack
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_plus_offset/$entry
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_plus_offset/$exit
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_plus_offset/sum_rename_req
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_base_plus_offset/sum_rename_ack
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_word_addrgen/$entry
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_word_addrgen/$exit
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_word_addrgen/root_register_req
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_word_addrgen/root_register_ack
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Sample/$entry
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Sample/word_access_start/$entry
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Sample/word_access_start/word_0/$entry
      -- CP-element group 661: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Sample/word_access_start/word_0/rr
      -- 
    ack_9261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 661_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4177_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(661)); -- 
    rr_9294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(661), ack => ptr_deref_4181_load_0_req_0); -- 
    -- CP-element group 662:  transition  input  bypass 
    -- CP-element group 662: predecessors 
    -- CP-element group 662: 	661 
    -- CP-element group 662: successors 
    -- CP-element group 662:  members (5) 
      -- CP-element group 662: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_sample_completed_
      -- CP-element group 662: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Sample/$exit
      -- CP-element group 662: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Sample/word_access_start/$exit
      -- CP-element group 662: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Sample/word_access_start/word_0/$exit
      -- CP-element group 662: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Sample/word_access_start/word_0/ra
      -- 
    ra_9295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 662_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4181_load_0_ack_0, ack => zeropad3D_CP_2067_elements(662)); -- 
    -- CP-element group 663:  transition  input  bypass 
    -- CP-element group 663: predecessors 
    -- CP-element group 663: 	638 
    -- CP-element group 663: successors 
    -- CP-element group 663: 	670 
    -- CP-element group 663:  members (9) 
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_update_completed_
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/$exit
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/word_access_complete/$exit
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/word_access_complete/word_0/$exit
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/word_access_complete/word_0/ca
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/ptr_deref_4181_Merge/$entry
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/ptr_deref_4181_Merge/$exit
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/ptr_deref_4181_Merge/merge_req
      -- CP-element group 663: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4181_Update/ptr_deref_4181_Merge/merge_ack
      -- 
    ca_9306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 663_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4181_load_0_ack_1, ack => zeropad3D_CP_2067_elements(663)); -- 
    -- CP-element group 664:  transition  input  bypass 
    -- CP-element group 664: predecessors 
    -- CP-element group 664: 	655 
    -- CP-element group 664: successors 
    -- CP-element group 664:  members (3) 
      -- CP-element group 664: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_sample_completed_
      -- CP-element group 664: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_Sample/$exit
      -- CP-element group 664: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_Sample/ra
      -- 
    ra_9320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 664_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4195_inst_ack_0, ack => zeropad3D_CP_2067_elements(664)); -- 
    -- CP-element group 665:  transition  input  output  bypass 
    -- CP-element group 665: predecessors 
    -- CP-element group 665: 	638 
    -- CP-element group 665: successors 
    -- CP-element group 665: 	666 
    -- CP-element group 665:  members (16) 
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_update_completed_
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_Update/$exit
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/type_cast_4195_Update/ca
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_resized_1
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_scaled_1
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_computed_1
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_resize_1/$entry
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_resize_1/$exit
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_resize_1/index_resize_req
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_resize_1/index_resize_ack
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_scale_1/$entry
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_scale_1/$exit
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_scale_1/scale_rename_req
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_index_scale_1/scale_rename_ack
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_Sample/$entry
      -- CP-element group 665: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_Sample/req
      -- 
    ca_9325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 665_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4195_inst_ack_1, ack => zeropad3D_CP_2067_elements(665)); -- 
    req_9350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(665), ack => array_obj_ref_4201_index_offset_req_0); -- 
    -- CP-element group 666:  transition  input  bypass 
    -- CP-element group 666: predecessors 
    -- CP-element group 666: 	665 
    -- CP-element group 666: successors 
    -- CP-element group 666: 	673 
    -- CP-element group 666:  members (3) 
      -- CP-element group 666: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_sample_complete
      -- CP-element group 666: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_Sample/$exit
      -- CP-element group 666: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_Sample/ack
      -- 
    ack_9351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 666_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4201_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(666)); -- 
    -- CP-element group 667:  transition  input  output  bypass 
    -- CP-element group 667: predecessors 
    -- CP-element group 667: 	638 
    -- CP-element group 667: successors 
    -- CP-element group 667: 	668 
    -- CP-element group 667:  members (11) 
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_sample_start_
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_root_address_calculated
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_offset_calculated
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_Update/$exit
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_final_index_sum_regn_Update/ack
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_base_plus_offset/$entry
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_base_plus_offset/$exit
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_base_plus_offset/sum_rename_req
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/array_obj_ref_4201_base_plus_offset/sum_rename_ack
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_request/$entry
      -- CP-element group 667: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_request/req
      -- 
    ack_9356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 667_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4201_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(667)); -- 
    req_9365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(667), ack => addr_of_4202_final_reg_req_0); -- 
    -- CP-element group 668:  transition  input  bypass 
    -- CP-element group 668: predecessors 
    -- CP-element group 668: 	667 
    -- CP-element group 668: successors 
    -- CP-element group 668:  members (3) 
      -- CP-element group 668: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_sample_completed_
      -- CP-element group 668: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_request/$exit
      -- CP-element group 668: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_request/ack
      -- 
    ack_9366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 668_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4202_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(668)); -- 
    -- CP-element group 669:  fork  transition  input  bypass 
    -- CP-element group 669: predecessors 
    -- CP-element group 669: 	638 
    -- CP-element group 669: successors 
    -- CP-element group 669: 	670 
    -- CP-element group 669:  members (19) 
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_update_completed_
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_complete/$exit
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/addr_of_4202_complete/ack
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_address_calculated
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_word_address_calculated
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_root_address_calculated
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_address_resized
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_addr_resize/$entry
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_addr_resize/$exit
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_addr_resize/base_resize_req
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_addr_resize/base_resize_ack
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_plus_offset/$entry
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_plus_offset/$exit
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_plus_offset/sum_rename_req
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_base_plus_offset/sum_rename_ack
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_word_addrgen/$entry
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_word_addrgen/$exit
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_word_addrgen/root_register_req
      -- CP-element group 669: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_word_addrgen/root_register_ack
      -- 
    ack_9371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 669_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4202_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(669)); -- 
    -- CP-element group 670:  join  transition  output  bypass 
    -- CP-element group 670: predecessors 
    -- CP-element group 670: 	663 
    -- CP-element group 670: 	669 
    -- CP-element group 670: successors 
    -- CP-element group 670: 	671 
    -- CP-element group 670:  members (9) 
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_sample_start_
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/$entry
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/ptr_deref_4205_Split/$entry
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/ptr_deref_4205_Split/$exit
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/ptr_deref_4205_Split/split_req
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/ptr_deref_4205_Split/split_ack
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/word_access_start/$entry
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/word_access_start/word_0/$entry
      -- CP-element group 670: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/word_access_start/word_0/rr
      -- 
    rr_9409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(670), ack => ptr_deref_4205_store_0_req_0); -- 
    zeropad3D_cp_element_group_670: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_670"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(663) & zeropad3D_CP_2067_elements(669);
      gj_zeropad3D_cp_element_group_670 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(670), clk => clk, reset => reset); --
    end block;
    -- CP-element group 671:  transition  input  bypass 
    -- CP-element group 671: predecessors 
    -- CP-element group 671: 	670 
    -- CP-element group 671: successors 
    -- CP-element group 671:  members (5) 
      -- CP-element group 671: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_sample_completed_
      -- CP-element group 671: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/$exit
      -- CP-element group 671: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/word_access_start/$exit
      -- CP-element group 671: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/word_access_start/word_0/$exit
      -- CP-element group 671: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Sample/word_access_start/word_0/ra
      -- 
    ra_9410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 671_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4205_store_0_ack_0, ack => zeropad3D_CP_2067_elements(671)); -- 
    -- CP-element group 672:  transition  input  bypass 
    -- CP-element group 672: predecessors 
    -- CP-element group 672: 	638 
    -- CP-element group 672: successors 
    -- CP-element group 672: 	673 
    -- CP-element group 672:  members (5) 
      -- CP-element group 672: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_update_completed_
      -- CP-element group 672: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Update/$exit
      -- CP-element group 672: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Update/word_access_complete/$exit
      -- CP-element group 672: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Update/word_access_complete/word_0/$exit
      -- CP-element group 672: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/ptr_deref_4205_Update/word_access_complete/word_0/ca
      -- 
    ca_9421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 672_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4205_store_0_ack_1, ack => zeropad3D_CP_2067_elements(672)); -- 
    -- CP-element group 673:  join  transition  place  bypass 
    -- CP-element group 673: predecessors 
    -- CP-element group 673: 	658 
    -- CP-element group 673: 	666 
    -- CP-element group 673: 	672 
    -- CP-element group 673: successors 
    -- CP-element group 673: 	1165 
    -- CP-element group 673:  members (5) 
      -- CP-element group 673: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207__exit__
      -- CP-element group 673: 	 branch_block_stmt_655/ifx_xelse1387_ifx_xend1435
      -- CP-element group 673: 	 branch_block_stmt_655/assign_stmt_4107_to_assign_stmt_4207/$exit
      -- CP-element group 673: 	 branch_block_stmt_655/ifx_xelse1387_ifx_xend1435_PhiReq/$entry
      -- CP-element group 673: 	 branch_block_stmt_655/ifx_xelse1387_ifx_xend1435_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_673: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_673"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(658) & zeropad3D_CP_2067_elements(666) & zeropad3D_CP_2067_elements(672);
      gj_zeropad3D_cp_element_group_673 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(673), clk => clk, reset => reset); --
    end block;
    -- CP-element group 674:  transition  input  bypass 
    -- CP-element group 674: predecessors 
    -- CP-element group 674: 	1165 
    -- CP-element group 674: successors 
    -- CP-element group 674:  members (3) 
      -- CP-element group 674: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_sample_completed_
      -- CP-element group 674: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_Sample/$exit
      -- CP-element group 674: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_Sample/ra
      -- 
    ra_9433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 674_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4213_inst_ack_0, ack => zeropad3D_CP_2067_elements(674)); -- 
    -- CP-element group 675:  branch  transition  place  input  output  bypass 
    -- CP-element group 675: predecessors 
    -- CP-element group 675: 	1165 
    -- CP-element group 675: successors 
    -- CP-element group 675: 	676 
    -- CP-element group 675: 	677 
    -- CP-element group 675:  members (13) 
      -- CP-element group 675: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227__exit__
      -- CP-element group 675: 	 branch_block_stmt_655/if_stmt_4228__entry__
      -- CP-element group 675: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/$exit
      -- CP-element group 675: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_update_completed_
      -- CP-element group 675: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_Update/$exit
      -- CP-element group 675: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_Update/ca
      -- CP-element group 675: 	 branch_block_stmt_655/if_stmt_4228_dead_link/$entry
      -- CP-element group 675: 	 branch_block_stmt_655/if_stmt_4228_eval_test/$entry
      -- CP-element group 675: 	 branch_block_stmt_655/if_stmt_4228_eval_test/$exit
      -- CP-element group 675: 	 branch_block_stmt_655/if_stmt_4228_eval_test/branch_req
      -- CP-element group 675: 	 branch_block_stmt_655/R_cmp1443_4229_place
      -- CP-element group 675: 	 branch_block_stmt_655/if_stmt_4228_if_link/$entry
      -- CP-element group 675: 	 branch_block_stmt_655/if_stmt_4228_else_link/$entry
      -- 
    ca_9438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 675_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4213_inst_ack_1, ack => zeropad3D_CP_2067_elements(675)); -- 
    branch_req_9446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(675), ack => if_stmt_4228_branch_req_0); -- 
    -- CP-element group 676:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 676: predecessors 
    -- CP-element group 676: 	675 
    -- CP-element group 676: successors 
    -- CP-element group 676: 	1174 
    -- CP-element group 676: 	1175 
    -- CP-element group 676: 	1177 
    -- CP-element group 676: 	1178 
    -- CP-element group 676: 	1180 
    -- CP-element group 676: 	1181 
    -- CP-element group 676:  members (40) 
      -- CP-element group 676: 	 branch_block_stmt_655/assign_stmt_4240__entry__
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486
      -- CP-element group 676: 	 branch_block_stmt_655/assign_stmt_4240__exit__
      -- CP-element group 676: 	 branch_block_stmt_655/merge_stmt_4234__exit__
      -- CP-element group 676: 	 branch_block_stmt_655/if_stmt_4228_if_link/$exit
      -- CP-element group 676: 	 branch_block_stmt_655/if_stmt_4228_if_link/if_choice_transition
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xend1435_ifx_xthen1445
      -- CP-element group 676: 	 branch_block_stmt_655/assign_stmt_4240/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/assign_stmt_4240/$exit
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xend1435_ifx_xthen1445_PhiReq/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xend1435_ifx_xthen1445_PhiReq/$exit
      -- CP-element group 676: 	 branch_block_stmt_655/merge_stmt_4234_PhiReqMerge
      -- CP-element group 676: 	 branch_block_stmt_655/merge_stmt_4234_PhiAck/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/merge_stmt_4234_PhiAck/$exit
      -- CP-element group 676: 	 branch_block_stmt_655/merge_stmt_4234_PhiAck/dummy
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/Sample/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/Sample/rr
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/Update/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/Update/cr
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/Sample/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/Sample/rr
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/Update/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/Update/cr
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/Sample/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/Sample/rr
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/Update/$entry
      -- CP-element group 676: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/Update/cr
      -- 
    if_choice_transition_9451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 676_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4228_branch_ack_1, ack => zeropad3D_CP_2067_elements(676)); -- 
    rr_13485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(676), ack => type_cast_4325_inst_req_0); -- 
    cr_13490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(676), ack => type_cast_4325_inst_req_1); -- 
    rr_13508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(676), ack => type_cast_4332_inst_req_0); -- 
    cr_13513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(676), ack => type_cast_4332_inst_req_1); -- 
    rr_13531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(676), ack => type_cast_4338_inst_req_0); -- 
    cr_13536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(676), ack => type_cast_4338_inst_req_1); -- 
    -- CP-element group 677:  fork  transition  place  input  output  bypass 
    -- CP-element group 677: predecessors 
    -- CP-element group 677: 	675 
    -- CP-element group 677: successors 
    -- CP-element group 677: 	678 
    -- CP-element group 677: 	679 
    -- CP-element group 677: 	680 
    -- CP-element group 677: 	681 
    -- CP-element group 677: 	683 
    -- CP-element group 677: 	686 
    -- CP-element group 677: 	688 
    -- CP-element group 677: 	689 
    -- CP-element group 677: 	690 
    -- CP-element group 677: 	692 
    -- CP-element group 677:  members (54) 
      -- CP-element group 677: 	 branch_block_stmt_655/merge_stmt_4242__exit__
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314__entry__
      -- CP-element group 677: 	 branch_block_stmt_655/if_stmt_4228_else_link/$exit
      -- CP-element group 677: 	 branch_block_stmt_655/if_stmt_4228_else_link/else_choice_transition
      -- CP-element group 677: 	 branch_block_stmt_655/ifx_xend1435_ifx_xelse1450
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_sample_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_update_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_Sample/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_Sample/rr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_Update/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_Update/cr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_sample_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_update_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_word_address_calculated
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_root_address_calculated
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Sample/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Sample/word_access_start/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Sample/word_access_start/word_0/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Sample/word_access_start/word_0/rr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/word_access_complete/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/word_access_complete/word_0/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/word_access_complete/word_0/cr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_update_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_Update/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_Update/cr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_update_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_Update/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_Update/cr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_update_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_Update/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_Update/cr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_sample_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_update_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_word_address_calculated
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_root_address_calculated
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Sample/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Sample/word_access_start/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Sample/word_access_start/word_0/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Sample/word_access_start/word_0/rr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/word_access_complete/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/word_access_complete/word_0/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/word_access_complete/word_0/cr
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_update_start_
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_Update/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_Update/cr
      -- CP-element group 677: 	 branch_block_stmt_655/ifx_xend1435_ifx_xelse1450_PhiReq/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/ifx_xend1435_ifx_xelse1450_PhiReq/$exit
      -- CP-element group 677: 	 branch_block_stmt_655/merge_stmt_4242_PhiReqMerge
      -- CP-element group 677: 	 branch_block_stmt_655/merge_stmt_4242_PhiAck/$entry
      -- CP-element group 677: 	 branch_block_stmt_655/merge_stmt_4242_PhiAck/$exit
      -- CP-element group 677: 	 branch_block_stmt_655/merge_stmt_4242_PhiAck/dummy
      -- 
    else_choice_transition_9455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 677_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4228_branch_ack_0, ack => zeropad3D_CP_2067_elements(677)); -- 
    rr_9471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => type_cast_4252_inst_req_0); -- 
    cr_9476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => type_cast_4252_inst_req_1); -- 
    rr_9493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => LOAD_col_high_4255_load_0_req_0); -- 
    cr_9504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => LOAD_col_high_4255_load_0_req_1); -- 
    cr_9523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => type_cast_4259_inst_req_1); -- 
    cr_9537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => type_cast_4279_inst_req_1); -- 
    cr_9551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => type_cast_4296_inst_req_1); -- 
    rr_9568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => LOAD_row_high_4299_load_0_req_0); -- 
    cr_9579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => LOAD_row_high_4299_load_0_req_1); -- 
    cr_9598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(677), ack => type_cast_4303_inst_req_1); -- 
    -- CP-element group 678:  transition  input  bypass 
    -- CP-element group 678: predecessors 
    -- CP-element group 678: 	677 
    -- CP-element group 678: successors 
    -- CP-element group 678:  members (3) 
      -- CP-element group 678: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_sample_completed_
      -- CP-element group 678: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_Sample/$exit
      -- CP-element group 678: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_Sample/ra
      -- 
    ra_9472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 678_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4252_inst_ack_0, ack => zeropad3D_CP_2067_elements(678)); -- 
    -- CP-element group 679:  transition  input  bypass 
    -- CP-element group 679: predecessors 
    -- CP-element group 679: 	677 
    -- CP-element group 679: successors 
    -- CP-element group 679: 	684 
    -- CP-element group 679:  members (3) 
      -- CP-element group 679: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_update_completed_
      -- CP-element group 679: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_Update/$exit
      -- CP-element group 679: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4252_Update/ca
      -- 
    ca_9477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 679_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4252_inst_ack_1, ack => zeropad3D_CP_2067_elements(679)); -- 
    -- CP-element group 680:  transition  input  bypass 
    -- CP-element group 680: predecessors 
    -- CP-element group 680: 	677 
    -- CP-element group 680: successors 
    -- CP-element group 680:  members (5) 
      -- CP-element group 680: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_sample_completed_
      -- CP-element group 680: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Sample/$exit
      -- CP-element group 680: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Sample/word_access_start/$exit
      -- CP-element group 680: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Sample/word_access_start/word_0/$exit
      -- CP-element group 680: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Sample/word_access_start/word_0/ra
      -- 
    ra_9494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 680_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4255_load_0_ack_0, ack => zeropad3D_CP_2067_elements(680)); -- 
    -- CP-element group 681:  transition  input  output  bypass 
    -- CP-element group 681: predecessors 
    -- CP-element group 681: 	677 
    -- CP-element group 681: successors 
    -- CP-element group 681: 	682 
    -- CP-element group 681:  members (12) 
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_update_completed_
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/$exit
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/word_access_complete/$exit
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/word_access_complete/word_0/$exit
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/word_access_complete/word_0/ca
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/LOAD_col_high_4255_Merge/$entry
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/LOAD_col_high_4255_Merge/$exit
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/LOAD_col_high_4255_Merge/merge_req
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_col_high_4255_Update/LOAD_col_high_4255_Merge/merge_ack
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_sample_start_
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_Sample/$entry
      -- CP-element group 681: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_Sample/rr
      -- 
    ca_9505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 681_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4255_load_0_ack_1, ack => zeropad3D_CP_2067_elements(681)); -- 
    rr_9518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(681), ack => type_cast_4259_inst_req_0); -- 
    -- CP-element group 682:  transition  input  bypass 
    -- CP-element group 682: predecessors 
    -- CP-element group 682: 	681 
    -- CP-element group 682: successors 
    -- CP-element group 682:  members (3) 
      -- CP-element group 682: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_sample_completed_
      -- CP-element group 682: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_Sample/$exit
      -- CP-element group 682: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_Sample/ra
      -- 
    ra_9519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 682_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4259_inst_ack_0, ack => zeropad3D_CP_2067_elements(682)); -- 
    -- CP-element group 683:  transition  input  bypass 
    -- CP-element group 683: predecessors 
    -- CP-element group 683: 	677 
    -- CP-element group 683: successors 
    -- CP-element group 683: 	684 
    -- CP-element group 683:  members (3) 
      -- CP-element group 683: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_update_completed_
      -- CP-element group 683: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_Update/$exit
      -- CP-element group 683: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4259_Update/ca
      -- 
    ca_9524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 683_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4259_inst_ack_1, ack => zeropad3D_CP_2067_elements(683)); -- 
    -- CP-element group 684:  join  transition  output  bypass 
    -- CP-element group 684: predecessors 
    -- CP-element group 684: 	679 
    -- CP-element group 684: 	683 
    -- CP-element group 684: successors 
    -- CP-element group 684: 	685 
    -- CP-element group 684:  members (3) 
      -- CP-element group 684: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_sample_start_
      -- CP-element group 684: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_Sample/$entry
      -- CP-element group 684: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_Sample/rr
      -- 
    rr_9532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(684), ack => type_cast_4279_inst_req_0); -- 
    zeropad3D_cp_element_group_684: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_684"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(679) & zeropad3D_CP_2067_elements(683);
      gj_zeropad3D_cp_element_group_684 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(684), clk => clk, reset => reset); --
    end block;
    -- CP-element group 685:  transition  input  bypass 
    -- CP-element group 685: predecessors 
    -- CP-element group 685: 	684 
    -- CP-element group 685: successors 
    -- CP-element group 685:  members (3) 
      -- CP-element group 685: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_sample_completed_
      -- CP-element group 685: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_Sample/$exit
      -- CP-element group 685: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_Sample/ra
      -- 
    ra_9533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 685_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4279_inst_ack_0, ack => zeropad3D_CP_2067_elements(685)); -- 
    -- CP-element group 686:  transition  input  output  bypass 
    -- CP-element group 686: predecessors 
    -- CP-element group 686: 	677 
    -- CP-element group 686: successors 
    -- CP-element group 686: 	687 
    -- CP-element group 686:  members (6) 
      -- CP-element group 686: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_update_completed_
      -- CP-element group 686: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_Update/$exit
      -- CP-element group 686: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4279_Update/ca
      -- CP-element group 686: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_sample_start_
      -- CP-element group 686: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_Sample/$entry
      -- CP-element group 686: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_Sample/rr
      -- 
    ca_9538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 686_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4279_inst_ack_1, ack => zeropad3D_CP_2067_elements(686)); -- 
    rr_9546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(686), ack => type_cast_4296_inst_req_0); -- 
    -- CP-element group 687:  transition  input  bypass 
    -- CP-element group 687: predecessors 
    -- CP-element group 687: 	686 
    -- CP-element group 687: successors 
    -- CP-element group 687:  members (3) 
      -- CP-element group 687: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_sample_completed_
      -- CP-element group 687: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_Sample/$exit
      -- CP-element group 687: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_Sample/ra
      -- 
    ra_9547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 687_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4296_inst_ack_0, ack => zeropad3D_CP_2067_elements(687)); -- 
    -- CP-element group 688:  transition  input  bypass 
    -- CP-element group 688: predecessors 
    -- CP-element group 688: 	677 
    -- CP-element group 688: successors 
    -- CP-element group 688: 	693 
    -- CP-element group 688:  members (3) 
      -- CP-element group 688: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_update_completed_
      -- CP-element group 688: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_Update/$exit
      -- CP-element group 688: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4296_Update/ca
      -- 
    ca_9552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 688_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4296_inst_ack_1, ack => zeropad3D_CP_2067_elements(688)); -- 
    -- CP-element group 689:  transition  input  bypass 
    -- CP-element group 689: predecessors 
    -- CP-element group 689: 	677 
    -- CP-element group 689: successors 
    -- CP-element group 689:  members (5) 
      -- CP-element group 689: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_sample_completed_
      -- CP-element group 689: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Sample/$exit
      -- CP-element group 689: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Sample/word_access_start/$exit
      -- CP-element group 689: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Sample/word_access_start/word_0/$exit
      -- CP-element group 689: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Sample/word_access_start/word_0/ra
      -- 
    ra_9569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 689_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4299_load_0_ack_0, ack => zeropad3D_CP_2067_elements(689)); -- 
    -- CP-element group 690:  transition  input  output  bypass 
    -- CP-element group 690: predecessors 
    -- CP-element group 690: 	677 
    -- CP-element group 690: successors 
    -- CP-element group 690: 	691 
    -- CP-element group 690:  members (12) 
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_update_completed_
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/$exit
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/word_access_complete/$exit
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/word_access_complete/word_0/$exit
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/word_access_complete/word_0/ca
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/LOAD_row_high_4299_Merge/$entry
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/LOAD_row_high_4299_Merge/$exit
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/LOAD_row_high_4299_Merge/merge_req
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/LOAD_row_high_4299_Update/LOAD_row_high_4299_Merge/merge_ack
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_sample_start_
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_Sample/$entry
      -- CP-element group 690: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_Sample/rr
      -- 
    ca_9580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 690_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4299_load_0_ack_1, ack => zeropad3D_CP_2067_elements(690)); -- 
    rr_9593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(690), ack => type_cast_4303_inst_req_0); -- 
    -- CP-element group 691:  transition  input  bypass 
    -- CP-element group 691: predecessors 
    -- CP-element group 691: 	690 
    -- CP-element group 691: successors 
    -- CP-element group 691:  members (3) 
      -- CP-element group 691: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_sample_completed_
      -- CP-element group 691: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_Sample/$exit
      -- CP-element group 691: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_Sample/ra
      -- 
    ra_9594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 691_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4303_inst_ack_0, ack => zeropad3D_CP_2067_elements(691)); -- 
    -- CP-element group 692:  transition  input  bypass 
    -- CP-element group 692: predecessors 
    -- CP-element group 692: 	677 
    -- CP-element group 692: successors 
    -- CP-element group 692: 	693 
    -- CP-element group 692:  members (3) 
      -- CP-element group 692: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_update_completed_
      -- CP-element group 692: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_Update/$exit
      -- CP-element group 692: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/type_cast_4303_Update/ca
      -- 
    ca_9599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 692_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4303_inst_ack_1, ack => zeropad3D_CP_2067_elements(692)); -- 
    -- CP-element group 693:  branch  join  transition  place  output  bypass 
    -- CP-element group 693: predecessors 
    -- CP-element group 693: 	688 
    -- CP-element group 693: 	692 
    -- CP-element group 693: successors 
    -- CP-element group 693: 	694 
    -- CP-element group 693: 	695 
    -- CP-element group 693:  members (10) 
      -- CP-element group 693: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314__exit__
      -- CP-element group 693: 	 branch_block_stmt_655/if_stmt_4315__entry__
      -- CP-element group 693: 	 branch_block_stmt_655/assign_stmt_4248_to_assign_stmt_4314/$exit
      -- CP-element group 693: 	 branch_block_stmt_655/if_stmt_4315_dead_link/$entry
      -- CP-element group 693: 	 branch_block_stmt_655/if_stmt_4315_eval_test/$entry
      -- CP-element group 693: 	 branch_block_stmt_655/if_stmt_4315_eval_test/$exit
      -- CP-element group 693: 	 branch_block_stmt_655/if_stmt_4315_eval_test/branch_req
      -- CP-element group 693: 	 branch_block_stmt_655/R_cmp1477_4316_place
      -- CP-element group 693: 	 branch_block_stmt_655/if_stmt_4315_if_link/$entry
      -- CP-element group 693: 	 branch_block_stmt_655/if_stmt_4315_else_link/$entry
      -- 
    branch_req_9607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(693), ack => if_stmt_4315_branch_req_0); -- 
    zeropad3D_cp_element_group_693: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_693"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(688) & zeropad3D_CP_2067_elements(692);
      gj_zeropad3D_cp_element_group_693 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(693), clk => clk, reset => reset); --
    end block;
    -- CP-element group 694:  fork  transition  place  input  output  bypass 
    -- CP-element group 694: predecessors 
    -- CP-element group 694: 	693 
    -- CP-element group 694: successors 
    -- CP-element group 694: 	1189 
    -- CP-element group 694: 	1190 
    -- CP-element group 694: 	1192 
    -- CP-element group 694: 	1193 
    -- CP-element group 694: 	1195 
    -- CP-element group 694: 	1196 
    -- CP-element group 694:  members (28) 
      -- CP-element group 694: 	 branch_block_stmt_655/if_stmt_4315_if_link/$exit
      -- CP-element group 694: 	 branch_block_stmt_655/if_stmt_4315_if_link/if_choice_transition
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/Sample/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/Sample/rr
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/Update/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/Update/cr
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/Sample/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/Sample/rr
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/Update/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/Update/cr
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Sample/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Sample/rr
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Update/$entry
      -- CP-element group 694: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Update/cr
      -- 
    if_choice_transition_9612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 694_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4315_branch_ack_1, ack => zeropad3D_CP_2067_elements(694)); -- 
    rr_13564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(694), ack => type_cast_4347_inst_req_0); -- 
    cr_13569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(694), ack => type_cast_4347_inst_req_1); -- 
    rr_13587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(694), ack => type_cast_4351_inst_req_0); -- 
    cr_13592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(694), ack => type_cast_4351_inst_req_1); -- 
    rr_13610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(694), ack => type_cast_4355_inst_req_0); -- 
    cr_13615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(694), ack => type_cast_4355_inst_req_1); -- 
    -- CP-element group 695:  fork  transition  place  input  output  bypass 
    -- CP-element group 695: predecessors 
    -- CP-element group 695: 	693 
    -- CP-element group 695: successors 
    -- CP-element group 695: 	1166 
    -- CP-element group 695: 	1167 
    -- CP-element group 695: 	1168 
    -- CP-element group 695: 	1170 
    -- CP-element group 695: 	1171 
    -- CP-element group 695:  members (22) 
      -- CP-element group 695: 	 branch_block_stmt_655/if_stmt_4315_else_link/$exit
      -- CP-element group 695: 	 branch_block_stmt_655/if_stmt_4315_else_link/else_choice_transition
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4322/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/Sample/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/Sample/rr
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/Update/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/Update/cr
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/Sample/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/Sample/rr
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/Update/$entry
      -- CP-element group 695: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/Update/cr
      -- 
    else_choice_transition_9616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 695_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4315_branch_ack_0, ack => zeropad3D_CP_2067_elements(695)); -- 
    rr_13436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(695), ack => type_cast_4334_inst_req_0); -- 
    cr_13441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(695), ack => type_cast_4334_inst_req_1); -- 
    rr_13459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(695), ack => type_cast_4340_inst_req_0); -- 
    cr_13464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(695), ack => type_cast_4340_inst_req_1); -- 
    -- CP-element group 696:  transition  input  bypass 
    -- CP-element group 696: predecessors 
    -- CP-element group 696: 	1202 
    -- CP-element group 696: successors 
    -- CP-element group 696:  members (3) 
      -- CP-element group 696: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_sample_completed_
      -- CP-element group 696: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_Sample/$exit
      -- CP-element group 696: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_Sample/ra
      -- 
    ra_9630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 696_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4359_inst_ack_0, ack => zeropad3D_CP_2067_elements(696)); -- 
    -- CP-element group 697:  transition  input  bypass 
    -- CP-element group 697: predecessors 
    -- CP-element group 697: 	1202 
    -- CP-element group 697: successors 
    -- CP-element group 697: 	718 
    -- CP-element group 697:  members (3) 
      -- CP-element group 697: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_update_completed_
      -- CP-element group 697: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_Update/$exit
      -- CP-element group 697: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_Update/ca
      -- 
    ca_9635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 697_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4359_inst_ack_1, ack => zeropad3D_CP_2067_elements(697)); -- 
    -- CP-element group 698:  transition  input  bypass 
    -- CP-element group 698: predecessors 
    -- CP-element group 698: 	1202 
    -- CP-element group 698: successors 
    -- CP-element group 698:  members (3) 
      -- CP-element group 698: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_sample_completed_
      -- CP-element group 698: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_Sample/$exit
      -- CP-element group 698: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_Sample/ra
      -- 
    ra_9644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 698_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4369_inst_ack_0, ack => zeropad3D_CP_2067_elements(698)); -- 
    -- CP-element group 699:  transition  input  bypass 
    -- CP-element group 699: predecessors 
    -- CP-element group 699: 	1202 
    -- CP-element group 699: successors 
    -- CP-element group 699: 	718 
    -- CP-element group 699:  members (3) 
      -- CP-element group 699: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_update_completed_
      -- CP-element group 699: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_Update/$exit
      -- CP-element group 699: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_Update/ca
      -- 
    ca_9649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 699_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4369_inst_ack_1, ack => zeropad3D_CP_2067_elements(699)); -- 
    -- CP-element group 700:  transition  input  bypass 
    -- CP-element group 700: predecessors 
    -- CP-element group 700: 	1202 
    -- CP-element group 700: successors 
    -- CP-element group 700:  members (5) 
      -- CP-element group 700: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_sample_completed_
      -- CP-element group 700: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Sample/$exit
      -- CP-element group 700: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Sample/word_access_start/$exit
      -- CP-element group 700: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Sample/word_access_start/word_0/$exit
      -- CP-element group 700: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Sample/word_access_start/word_0/ra
      -- 
    ra_9666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 700_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4384_load_0_ack_0, ack => zeropad3D_CP_2067_elements(700)); -- 
    -- CP-element group 701:  transition  input  output  bypass 
    -- CP-element group 701: predecessors 
    -- CP-element group 701: 	1202 
    -- CP-element group 701: successors 
    -- CP-element group 701: 	714 
    -- CP-element group 701:  members (12) 
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_update_completed_
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/$exit
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/word_access_complete/$exit
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/word_access_complete/word_0/$exit
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/word_access_complete/word_0/ca
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/LOAD_pad_4384_Merge/$entry
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/LOAD_pad_4384_Merge/$exit
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/LOAD_pad_4384_Merge/merge_req
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/LOAD_pad_4384_Merge/merge_ack
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_sample_start_
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_Sample/$entry
      -- CP-element group 701: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_Sample/rr
      -- 
    ca_9677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 701_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4384_load_0_ack_1, ack => zeropad3D_CP_2067_elements(701)); -- 
    rr_9831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(701), ack => type_cast_4414_inst_req_0); -- 
    -- CP-element group 702:  transition  input  bypass 
    -- CP-element group 702: predecessors 
    -- CP-element group 702: 	1202 
    -- CP-element group 702: successors 
    -- CP-element group 702:  members (5) 
      -- CP-element group 702: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_sample_completed_
      -- CP-element group 702: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Sample/$exit
      -- CP-element group 702: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Sample/word_access_start/$exit
      -- CP-element group 702: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Sample/word_access_start/word_0/$exit
      -- CP-element group 702: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Sample/word_access_start/word_0/ra
      -- 
    ra_9699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 702_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4387_load_0_ack_0, ack => zeropad3D_CP_2067_elements(702)); -- 
    -- CP-element group 703:  transition  input  output  bypass 
    -- CP-element group 703: predecessors 
    -- CP-element group 703: 	1202 
    -- CP-element group 703: successors 
    -- CP-element group 703: 	708 
    -- CP-element group 703:  members (12) 
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_update_completed_
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/$exit
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/word_access_complete/$exit
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/word_access_complete/word_0/$exit
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/word_access_complete/word_0/ca
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/LOAD_depth_high_4387_Merge/$entry
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/LOAD_depth_high_4387_Merge/$exit
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/LOAD_depth_high_4387_Merge/merge_req
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/LOAD_depth_high_4387_Merge/merge_ack
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_sample_start_
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_Sample/$entry
      -- CP-element group 703: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_Sample/rr
      -- 
    ca_9710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 703_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4387_load_0_ack_1, ack => zeropad3D_CP_2067_elements(703)); -- 
    rr_9789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(703), ack => type_cast_4397_inst_req_0); -- 
    -- CP-element group 704:  transition  input  bypass 
    -- CP-element group 704: predecessors 
    -- CP-element group 704: 	1202 
    -- CP-element group 704: successors 
    -- CP-element group 704:  members (5) 
      -- CP-element group 704: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_sample_completed_
      -- CP-element group 704: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Sample/$exit
      -- CP-element group 704: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Sample/word_access_start/$exit
      -- CP-element group 704: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Sample/word_access_start/word_0/$exit
      -- CP-element group 704: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Sample/word_access_start/word_0/ra
      -- 
    ra_9732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 704_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_4390_load_0_ack_0, ack => zeropad3D_CP_2067_elements(704)); -- 
    -- CP-element group 705:  fork  transition  input  output  bypass 
    -- CP-element group 705: predecessors 
    -- CP-element group 705: 	1202 
    -- CP-element group 705: successors 
    -- CP-element group 705: 	710 
    -- CP-element group 705: 	716 
    -- CP-element group 705:  members (15) 
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_update_completed_
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/$exit
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/word_access_complete/$exit
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/word_access_complete/word_0/$exit
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/word_access_complete/word_0/ca
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/LOAD_out_depth_high_4390_Merge/$entry
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/LOAD_out_depth_high_4390_Merge/$exit
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/LOAD_out_depth_high_4390_Merge/merge_req
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/LOAD_out_depth_high_4390_Merge/merge_ack
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_sample_start_
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_Sample/$entry
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_Sample/rr
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_sample_start_
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_Sample/$entry
      -- CP-element group 705: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_Sample/rr
      -- 
    ca_9743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 705_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_depth_high_4390_load_0_ack_1, ack => zeropad3D_CP_2067_elements(705)); -- 
    rr_9803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(705), ack => type_cast_4401_inst_req_0); -- 
    rr_9845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(705), ack => type_cast_4418_inst_req_0); -- 
    -- CP-element group 706:  transition  input  bypass 
    -- CP-element group 706: predecessors 
    -- CP-element group 706: 	1202 
    -- CP-element group 706: successors 
    -- CP-element group 706:  members (5) 
      -- CP-element group 706: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_sample_completed_
      -- CP-element group 706: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Sample/$exit
      -- CP-element group 706: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Sample/word_access_start/$exit
      -- CP-element group 706: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Sample/word_access_start/word_0/$exit
      -- CP-element group 706: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Sample/word_access_start/word_0/ra
      -- 
    ra_9765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 706_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_4393_load_0_ack_0, ack => zeropad3D_CP_2067_elements(706)); -- 
    -- CP-element group 707:  transition  input  output  bypass 
    -- CP-element group 707: predecessors 
    -- CP-element group 707: 	1202 
    -- CP-element group 707: successors 
    -- CP-element group 707: 	712 
    -- CP-element group 707:  members (12) 
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_update_completed_
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/$exit
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/word_access_complete/$exit
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/word_access_complete/word_0/$exit
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/word_access_complete/word_0/ca
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/LOAD_out_col_high_4393_Merge/$entry
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/LOAD_out_col_high_4393_Merge/$exit
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/LOAD_out_col_high_4393_Merge/merge_req
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/LOAD_out_col_high_4393_Merge/merge_ack
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_sample_start_
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_Sample/$entry
      -- CP-element group 707: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_Sample/rr
      -- 
    ca_9776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 707_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_out_col_high_4393_load_0_ack_1, ack => zeropad3D_CP_2067_elements(707)); -- 
    rr_9817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(707), ack => type_cast_4405_inst_req_0); -- 
    -- CP-element group 708:  transition  input  bypass 
    -- CP-element group 708: predecessors 
    -- CP-element group 708: 	703 
    -- CP-element group 708: successors 
    -- CP-element group 708:  members (3) 
      -- CP-element group 708: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_sample_completed_
      -- CP-element group 708: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_Sample/$exit
      -- CP-element group 708: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_Sample/ra
      -- 
    ra_9790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 708_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4397_inst_ack_0, ack => zeropad3D_CP_2067_elements(708)); -- 
    -- CP-element group 709:  transition  input  bypass 
    -- CP-element group 709: predecessors 
    -- CP-element group 709: 	1202 
    -- CP-element group 709: successors 
    -- CP-element group 709: 	718 
    -- CP-element group 709:  members (3) 
      -- CP-element group 709: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_update_completed_
      -- CP-element group 709: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_Update/$exit
      -- CP-element group 709: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_Update/ca
      -- 
    ca_9795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 709_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4397_inst_ack_1, ack => zeropad3D_CP_2067_elements(709)); -- 
    -- CP-element group 710:  transition  input  bypass 
    -- CP-element group 710: predecessors 
    -- CP-element group 710: 	705 
    -- CP-element group 710: successors 
    -- CP-element group 710:  members (3) 
      -- CP-element group 710: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_sample_completed_
      -- CP-element group 710: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_Sample/$exit
      -- CP-element group 710: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_Sample/ra
      -- 
    ra_9804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 710_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4401_inst_ack_0, ack => zeropad3D_CP_2067_elements(710)); -- 
    -- CP-element group 711:  transition  input  bypass 
    -- CP-element group 711: predecessors 
    -- CP-element group 711: 	1202 
    -- CP-element group 711: successors 
    -- CP-element group 711: 	718 
    -- CP-element group 711:  members (3) 
      -- CP-element group 711: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_update_completed_
      -- CP-element group 711: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_Update/$exit
      -- CP-element group 711: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_Update/ca
      -- 
    ca_9809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 711_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4401_inst_ack_1, ack => zeropad3D_CP_2067_elements(711)); -- 
    -- CP-element group 712:  transition  input  bypass 
    -- CP-element group 712: predecessors 
    -- CP-element group 712: 	707 
    -- CP-element group 712: successors 
    -- CP-element group 712:  members (3) 
      -- CP-element group 712: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_sample_completed_
      -- CP-element group 712: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_Sample/$exit
      -- CP-element group 712: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_Sample/ra
      -- 
    ra_9818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 712_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4405_inst_ack_0, ack => zeropad3D_CP_2067_elements(712)); -- 
    -- CP-element group 713:  transition  input  bypass 
    -- CP-element group 713: predecessors 
    -- CP-element group 713: 	1202 
    -- CP-element group 713: successors 
    -- CP-element group 713: 	718 
    -- CP-element group 713:  members (3) 
      -- CP-element group 713: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_update_completed_
      -- CP-element group 713: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_Update/$exit
      -- CP-element group 713: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_Update/ca
      -- 
    ca_9823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 713_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4405_inst_ack_1, ack => zeropad3D_CP_2067_elements(713)); -- 
    -- CP-element group 714:  transition  input  bypass 
    -- CP-element group 714: predecessors 
    -- CP-element group 714: 	701 
    -- CP-element group 714: successors 
    -- CP-element group 714:  members (3) 
      -- CP-element group 714: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_sample_completed_
      -- CP-element group 714: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_Sample/$exit
      -- CP-element group 714: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_Sample/ra
      -- 
    ra_9832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 714_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4414_inst_ack_0, ack => zeropad3D_CP_2067_elements(714)); -- 
    -- CP-element group 715:  transition  input  bypass 
    -- CP-element group 715: predecessors 
    -- CP-element group 715: 	1202 
    -- CP-element group 715: successors 
    -- CP-element group 715: 	718 
    -- CP-element group 715:  members (3) 
      -- CP-element group 715: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_update_completed_
      -- CP-element group 715: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_Update/$exit
      -- CP-element group 715: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_Update/ca
      -- 
    ca_9837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 715_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4414_inst_ack_1, ack => zeropad3D_CP_2067_elements(715)); -- 
    -- CP-element group 716:  transition  input  bypass 
    -- CP-element group 716: predecessors 
    -- CP-element group 716: 	705 
    -- CP-element group 716: successors 
    -- CP-element group 716:  members (3) 
      -- CP-element group 716: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_sample_completed_
      -- CP-element group 716: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_Sample/$exit
      -- CP-element group 716: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_Sample/ra
      -- 
    ra_9846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 716_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4418_inst_ack_0, ack => zeropad3D_CP_2067_elements(716)); -- 
    -- CP-element group 717:  transition  input  bypass 
    -- CP-element group 717: predecessors 
    -- CP-element group 717: 	1202 
    -- CP-element group 717: successors 
    -- CP-element group 717: 	718 
    -- CP-element group 717:  members (3) 
      -- CP-element group 717: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_update_completed_
      -- CP-element group 717: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_Update/$exit
      -- CP-element group 717: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_Update/ca
      -- 
    ca_9851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 717_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4418_inst_ack_1, ack => zeropad3D_CP_2067_elements(717)); -- 
    -- CP-element group 718:  join  fork  transition  place  output  bypass 
    -- CP-element group 718: predecessors 
    -- CP-element group 718: 	697 
    -- CP-element group 718: 	699 
    -- CP-element group 718: 	709 
    -- CP-element group 718: 	711 
    -- CP-element group 718: 	713 
    -- CP-element group 718: 	715 
    -- CP-element group 718: 	717 
    -- CP-element group 718: successors 
    -- CP-element group 718: 	1213 
    -- CP-element group 718: 	1214 
    -- CP-element group 718: 	1215 
    -- CP-element group 718: 	1217 
    -- CP-element group 718: 	1218 
    -- CP-element group 718:  members (22) 
      -- CP-element group 718: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460__exit__
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552
      -- CP-element group 718: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/$exit
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4463/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/Sample/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/Sample/rr
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/Update/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/Update/cr
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/Sample/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/Sample/rr
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/Update/$entry
      -- CP-element group 718: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/Update/cr
      -- 
    rr_13723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(718), ack => type_cast_4473_inst_req_0); -- 
    cr_13728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(718), ack => type_cast_4473_inst_req_1); -- 
    rr_13746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(718), ack => type_cast_4479_inst_req_0); -- 
    cr_13751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(718), ack => type_cast_4479_inst_req_1); -- 
    zeropad3D_cp_element_group_718: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_718"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(697) & zeropad3D_CP_2067_elements(699) & zeropad3D_CP_2067_elements(709) & zeropad3D_CP_2067_elements(711) & zeropad3D_CP_2067_elements(713) & zeropad3D_CP_2067_elements(715) & zeropad3D_CP_2067_elements(717);
      gj_zeropad3D_cp_element_group_718 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(718), clk => clk, reset => reset); --
    end block;
    -- CP-element group 719:  transition  input  bypass 
    -- CP-element group 719: predecessors 
    -- CP-element group 719: 	1225 
    -- CP-element group 719: successors 
    -- CP-element group 719:  members (3) 
      -- CP-element group 719: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_sample_completed_
      -- CP-element group 719: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_Sample/$exit
      -- CP-element group 719: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_Sample/ra
      -- 
    ra_9863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 719_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4486_inst_ack_0, ack => zeropad3D_CP_2067_elements(719)); -- 
    -- CP-element group 720:  branch  transition  place  input  output  bypass 
    -- CP-element group 720: predecessors 
    -- CP-element group 720: 	1225 
    -- CP-element group 720: successors 
    -- CP-element group 720: 	721 
    -- CP-element group 720: 	722 
    -- CP-element group 720:  members (13) 
      -- CP-element group 720: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494__exit__
      -- CP-element group 720: 	 branch_block_stmt_655/if_stmt_4495__entry__
      -- CP-element group 720: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/$exit
      -- CP-element group 720: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_update_completed_
      -- CP-element group 720: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_Update/$exit
      -- CP-element group 720: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_Update/ca
      -- CP-element group 720: 	 branch_block_stmt_655/if_stmt_4495_dead_link/$entry
      -- CP-element group 720: 	 branch_block_stmt_655/if_stmt_4495_eval_test/$entry
      -- CP-element group 720: 	 branch_block_stmt_655/if_stmt_4495_eval_test/$exit
      -- CP-element group 720: 	 branch_block_stmt_655/if_stmt_4495_eval_test/branch_req
      -- CP-element group 720: 	 branch_block_stmt_655/R_cmp1557_4496_place
      -- CP-element group 720: 	 branch_block_stmt_655/if_stmt_4495_if_link/$entry
      -- CP-element group 720: 	 branch_block_stmt_655/if_stmt_4495_else_link/$entry
      -- 
    ca_9868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 720_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4486_inst_ack_1, ack => zeropad3D_CP_2067_elements(720)); -- 
    branch_req_9876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(720), ack => if_stmt_4495_branch_req_0); -- 
    -- CP-element group 721:  transition  place  input  bypass 
    -- CP-element group 721: predecessors 
    -- CP-element group 721: 	720 
    -- CP-element group 721: successors 
    -- CP-element group 721: 	1226 
    -- CP-element group 721:  members (5) 
      -- CP-element group 721: 	 branch_block_stmt_655/if_stmt_4495_if_link/$exit
      -- CP-element group 721: 	 branch_block_stmt_655/if_stmt_4495_if_link/if_choice_transition
      -- CP-element group 721: 	 branch_block_stmt_655/whilex_xbody1552_ifx_xthen1586
      -- CP-element group 721: 	 branch_block_stmt_655/whilex_xbody1552_ifx_xthen1586_PhiReq/$entry
      -- CP-element group 721: 	 branch_block_stmt_655/whilex_xbody1552_ifx_xthen1586_PhiReq/$exit
      -- 
    if_choice_transition_9881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 721_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4495_branch_ack_1, ack => zeropad3D_CP_2067_elements(721)); -- 
    -- CP-element group 722:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 722: predecessors 
    -- CP-element group 722: 	720 
    -- CP-element group 722: successors 
    -- CP-element group 722: 	723 
    -- CP-element group 722: 	724 
    -- CP-element group 722: 	726 
    -- CP-element group 722:  members (27) 
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520__entry__
      -- CP-element group 722: 	 branch_block_stmt_655/merge_stmt_4501__exit__
      -- CP-element group 722: 	 branch_block_stmt_655/if_stmt_4495_else_link/$exit
      -- CP-element group 722: 	 branch_block_stmt_655/if_stmt_4495_else_link/else_choice_transition
      -- CP-element group 722: 	 branch_block_stmt_655/whilex_xbody1552_lorx_xlhsx_xfalse1559
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_sample_start_
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_update_start_
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_word_address_calculated
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_root_address_calculated
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Sample/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Sample/word_access_start/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Sample/word_access_start/word_0/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Sample/word_access_start/word_0/rr
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/word_access_complete/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/word_access_complete/word_0/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/word_access_complete/word_0/cr
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_update_start_
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_655/whilex_xbody1552_lorx_xlhsx_xfalse1559_PhiReq/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/whilex_xbody1552_lorx_xlhsx_xfalse1559_PhiReq/$exit
      -- CP-element group 722: 	 branch_block_stmt_655/merge_stmt_4501_PhiReqMerge
      -- CP-element group 722: 	 branch_block_stmt_655/merge_stmt_4501_PhiAck/$entry
      -- CP-element group 722: 	 branch_block_stmt_655/merge_stmt_4501_PhiAck/$exit
      -- CP-element group 722: 	 branch_block_stmt_655/merge_stmt_4501_PhiAck/dummy
      -- 
    else_choice_transition_9885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 722_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4495_branch_ack_0, ack => zeropad3D_CP_2067_elements(722)); -- 
    rr_9906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(722), ack => LOAD_row_high_4503_load_0_req_0); -- 
    cr_9917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(722), ack => LOAD_row_high_4503_load_0_req_1); -- 
    cr_9936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(722), ack => type_cast_4507_inst_req_1); -- 
    -- CP-element group 723:  transition  input  bypass 
    -- CP-element group 723: predecessors 
    -- CP-element group 723: 	722 
    -- CP-element group 723: successors 
    -- CP-element group 723:  members (5) 
      -- CP-element group 723: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_sample_completed_
      -- CP-element group 723: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Sample/$exit
      -- CP-element group 723: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Sample/word_access_start/$exit
      -- CP-element group 723: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Sample/word_access_start/word_0/$exit
      -- CP-element group 723: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Sample/word_access_start/word_0/ra
      -- 
    ra_9907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 723_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4503_load_0_ack_0, ack => zeropad3D_CP_2067_elements(723)); -- 
    -- CP-element group 724:  transition  input  output  bypass 
    -- CP-element group 724: predecessors 
    -- CP-element group 724: 	722 
    -- CP-element group 724: successors 
    -- CP-element group 724: 	725 
    -- CP-element group 724:  members (12) 
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_update_completed_
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/$exit
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/word_access_complete/$exit
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/word_access_complete/word_0/$exit
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/word_access_complete/word_0/ca
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/LOAD_row_high_4503_Merge/$entry
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/LOAD_row_high_4503_Merge/$exit
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/LOAD_row_high_4503_Merge/merge_req
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/LOAD_row_high_4503_Update/LOAD_row_high_4503_Merge/merge_ack
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_sample_start_
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_Sample/$entry
      -- CP-element group 724: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_Sample/rr
      -- 
    ca_9918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 724_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4503_load_0_ack_1, ack => zeropad3D_CP_2067_elements(724)); -- 
    rr_9931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(724), ack => type_cast_4507_inst_req_0); -- 
    -- CP-element group 725:  transition  input  bypass 
    -- CP-element group 725: predecessors 
    -- CP-element group 725: 	724 
    -- CP-element group 725: successors 
    -- CP-element group 725:  members (3) 
      -- CP-element group 725: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_sample_completed_
      -- CP-element group 725: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_Sample/$exit
      -- CP-element group 725: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_Sample/ra
      -- 
    ra_9932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 725_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4507_inst_ack_0, ack => zeropad3D_CP_2067_elements(725)); -- 
    -- CP-element group 726:  branch  transition  place  input  output  bypass 
    -- CP-element group 726: predecessors 
    -- CP-element group 726: 	722 
    -- CP-element group 726: successors 
    -- CP-element group 726: 	727 
    -- CP-element group 726: 	728 
    -- CP-element group 726:  members (13) 
      -- CP-element group 726: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520__exit__
      -- CP-element group 726: 	 branch_block_stmt_655/if_stmt_4521__entry__
      -- CP-element group 726: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/$exit
      -- CP-element group 726: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_update_completed_
      -- CP-element group 726: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_Update/$exit
      -- CP-element group 726: 	 branch_block_stmt_655/assign_stmt_4504_to_assign_stmt_4520/type_cast_4507_Update/ca
      -- CP-element group 726: 	 branch_block_stmt_655/if_stmt_4521_dead_link/$entry
      -- CP-element group 726: 	 branch_block_stmt_655/if_stmt_4521_eval_test/$entry
      -- CP-element group 726: 	 branch_block_stmt_655/if_stmt_4521_eval_test/$exit
      -- CP-element group 726: 	 branch_block_stmt_655/if_stmt_4521_eval_test/branch_req
      -- CP-element group 726: 	 branch_block_stmt_655/R_cmp1567_4522_place
      -- CP-element group 726: 	 branch_block_stmt_655/if_stmt_4521_if_link/$entry
      -- CP-element group 726: 	 branch_block_stmt_655/if_stmt_4521_else_link/$entry
      -- 
    ca_9937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 726_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4507_inst_ack_1, ack => zeropad3D_CP_2067_elements(726)); -- 
    branch_req_9945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(726), ack => if_stmt_4521_branch_req_0); -- 
    -- CP-element group 727:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 727: predecessors 
    -- CP-element group 727: 	726 
    -- CP-element group 727: successors 
    -- CP-element group 727: 	729 
    -- CP-element group 727: 	730 
    -- CP-element group 727:  members (18) 
      -- CP-element group 727: 	 branch_block_stmt_655/merge_stmt_4527__exit__
      -- CP-element group 727: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539__entry__
      -- CP-element group 727: 	 branch_block_stmt_655/if_stmt_4521_if_link/$exit
      -- CP-element group 727: 	 branch_block_stmt_655/if_stmt_4521_if_link/if_choice_transition
      -- CP-element group 727: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1559_lorx_xlhsx_xfalse1569
      -- CP-element group 727: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/$entry
      -- CP-element group 727: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_sample_start_
      -- CP-element group 727: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_update_start_
      -- CP-element group 727: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_Sample/$entry
      -- CP-element group 727: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_Sample/rr
      -- CP-element group 727: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_Update/$entry
      -- CP-element group 727: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_Update/cr
      -- CP-element group 727: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1559_lorx_xlhsx_xfalse1569_PhiReq/$entry
      -- CP-element group 727: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1559_lorx_xlhsx_xfalse1569_PhiReq/$exit
      -- CP-element group 727: 	 branch_block_stmt_655/merge_stmt_4527_PhiReqMerge
      -- CP-element group 727: 	 branch_block_stmt_655/merge_stmt_4527_PhiAck/$entry
      -- CP-element group 727: 	 branch_block_stmt_655/merge_stmt_4527_PhiAck/$exit
      -- CP-element group 727: 	 branch_block_stmt_655/merge_stmt_4527_PhiAck/dummy
      -- 
    if_choice_transition_9950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 727_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4521_branch_ack_1, ack => zeropad3D_CP_2067_elements(727)); -- 
    rr_9967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(727), ack => type_cast_4531_inst_req_0); -- 
    cr_9972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(727), ack => type_cast_4531_inst_req_1); -- 
    -- CP-element group 728:  transition  place  input  bypass 
    -- CP-element group 728: predecessors 
    -- CP-element group 728: 	726 
    -- CP-element group 728: successors 
    -- CP-element group 728: 	1226 
    -- CP-element group 728:  members (5) 
      -- CP-element group 728: 	 branch_block_stmt_655/if_stmt_4521_else_link/$exit
      -- CP-element group 728: 	 branch_block_stmt_655/if_stmt_4521_else_link/else_choice_transition
      -- CP-element group 728: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1559_ifx_xthen1586
      -- CP-element group 728: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1559_ifx_xthen1586_PhiReq/$entry
      -- CP-element group 728: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1559_ifx_xthen1586_PhiReq/$exit
      -- 
    else_choice_transition_9954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 728_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4521_branch_ack_0, ack => zeropad3D_CP_2067_elements(728)); -- 
    -- CP-element group 729:  transition  input  bypass 
    -- CP-element group 729: predecessors 
    -- CP-element group 729: 	727 
    -- CP-element group 729: successors 
    -- CP-element group 729:  members (3) 
      -- CP-element group 729: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_sample_completed_
      -- CP-element group 729: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_Sample/$exit
      -- CP-element group 729: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_Sample/ra
      -- 
    ra_9968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 729_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4531_inst_ack_0, ack => zeropad3D_CP_2067_elements(729)); -- 
    -- CP-element group 730:  branch  transition  place  input  output  bypass 
    -- CP-element group 730: predecessors 
    -- CP-element group 730: 	727 
    -- CP-element group 730: successors 
    -- CP-element group 730: 	731 
    -- CP-element group 730: 	732 
    -- CP-element group 730:  members (13) 
      -- CP-element group 730: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539__exit__
      -- CP-element group 730: 	 branch_block_stmt_655/if_stmt_4540__entry__
      -- CP-element group 730: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/$exit
      -- CP-element group 730: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_update_completed_
      -- CP-element group 730: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_Update/$exit
      -- CP-element group 730: 	 branch_block_stmt_655/assign_stmt_4532_to_assign_stmt_4539/type_cast_4531_Update/ca
      -- CP-element group 730: 	 branch_block_stmt_655/if_stmt_4540_dead_link/$entry
      -- CP-element group 730: 	 branch_block_stmt_655/if_stmt_4540_eval_test/$entry
      -- CP-element group 730: 	 branch_block_stmt_655/if_stmt_4540_eval_test/$exit
      -- CP-element group 730: 	 branch_block_stmt_655/if_stmt_4540_eval_test/branch_req
      -- CP-element group 730: 	 branch_block_stmt_655/R_cmp1574_4541_place
      -- CP-element group 730: 	 branch_block_stmt_655/if_stmt_4540_if_link/$entry
      -- CP-element group 730: 	 branch_block_stmt_655/if_stmt_4540_else_link/$entry
      -- 
    ca_9973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 730_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4531_inst_ack_1, ack => zeropad3D_CP_2067_elements(730)); -- 
    branch_req_9981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(730), ack => if_stmt_4540_branch_req_0); -- 
    -- CP-element group 731:  transition  place  input  bypass 
    -- CP-element group 731: predecessors 
    -- CP-element group 731: 	730 
    -- CP-element group 731: successors 
    -- CP-element group 731: 	1226 
    -- CP-element group 731:  members (5) 
      -- CP-element group 731: 	 branch_block_stmt_655/if_stmt_4540_if_link/$exit
      -- CP-element group 731: 	 branch_block_stmt_655/if_stmt_4540_if_link/if_choice_transition
      -- CP-element group 731: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1569_ifx_xthen1586
      -- CP-element group 731: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1569_ifx_xthen1586_PhiReq/$entry
      -- CP-element group 731: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1569_ifx_xthen1586_PhiReq/$exit
      -- 
    if_choice_transition_9986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 731_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4540_branch_ack_1, ack => zeropad3D_CP_2067_elements(731)); -- 
    -- CP-element group 732:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 732: predecessors 
    -- CP-element group 732: 	730 
    -- CP-element group 732: successors 
    -- CP-element group 732: 	733 
    -- CP-element group 732: 	734 
    -- CP-element group 732: 	736 
    -- CP-element group 732:  members (27) 
      -- CP-element group 732: 	 branch_block_stmt_655/merge_stmt_4546__exit__
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565__entry__
      -- CP-element group 732: 	 branch_block_stmt_655/if_stmt_4540_else_link/$exit
      -- CP-element group 732: 	 branch_block_stmt_655/if_stmt_4540_else_link/else_choice_transition
      -- CP-element group 732: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1576
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_sample_start_
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_update_start_
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_word_address_calculated
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_root_address_calculated
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Sample/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Sample/word_access_start/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Sample/word_access_start/word_0/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Sample/word_access_start/word_0/rr
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/word_access_complete/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/word_access_complete/word_0/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/word_access_complete/word_0/cr
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_update_start_
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_Update/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_Update/cr
      -- CP-element group 732: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1576_PhiReq/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1576_PhiReq/$exit
      -- CP-element group 732: 	 branch_block_stmt_655/merge_stmt_4546_PhiReqMerge
      -- CP-element group 732: 	 branch_block_stmt_655/merge_stmt_4546_PhiAck/$entry
      -- CP-element group 732: 	 branch_block_stmt_655/merge_stmt_4546_PhiAck/$exit
      -- CP-element group 732: 	 branch_block_stmt_655/merge_stmt_4546_PhiAck/dummy
      -- 
    else_choice_transition_9990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 732_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4540_branch_ack_0, ack => zeropad3D_CP_2067_elements(732)); -- 
    rr_10011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(732), ack => LOAD_col_high_4548_load_0_req_0); -- 
    cr_10022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(732), ack => LOAD_col_high_4548_load_0_req_1); -- 
    cr_10041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(732), ack => type_cast_4552_inst_req_1); -- 
    -- CP-element group 733:  transition  input  bypass 
    -- CP-element group 733: predecessors 
    -- CP-element group 733: 	732 
    -- CP-element group 733: successors 
    -- CP-element group 733:  members (5) 
      -- CP-element group 733: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_sample_completed_
      -- CP-element group 733: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Sample/$exit
      -- CP-element group 733: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Sample/word_access_start/$exit
      -- CP-element group 733: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Sample/word_access_start/word_0/$exit
      -- CP-element group 733: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Sample/word_access_start/word_0/ra
      -- 
    ra_10012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 733_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4548_load_0_ack_0, ack => zeropad3D_CP_2067_elements(733)); -- 
    -- CP-element group 734:  transition  input  output  bypass 
    -- CP-element group 734: predecessors 
    -- CP-element group 734: 	732 
    -- CP-element group 734: successors 
    -- CP-element group 734: 	735 
    -- CP-element group 734:  members (12) 
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_update_completed_
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/$exit
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/word_access_complete/$exit
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/word_access_complete/word_0/$exit
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/word_access_complete/word_0/ca
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/LOAD_col_high_4548_Merge/$entry
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/LOAD_col_high_4548_Merge/$exit
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/LOAD_col_high_4548_Merge/merge_req
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/LOAD_col_high_4548_Update/LOAD_col_high_4548_Merge/merge_ack
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_sample_start_
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_Sample/$entry
      -- CP-element group 734: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_Sample/rr
      -- 
    ca_10023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 734_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4548_load_0_ack_1, ack => zeropad3D_CP_2067_elements(734)); -- 
    rr_10036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(734), ack => type_cast_4552_inst_req_0); -- 
    -- CP-element group 735:  transition  input  bypass 
    -- CP-element group 735: predecessors 
    -- CP-element group 735: 	734 
    -- CP-element group 735: successors 
    -- CP-element group 735:  members (3) 
      -- CP-element group 735: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_sample_completed_
      -- CP-element group 735: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_Sample/$exit
      -- CP-element group 735: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_Sample/ra
      -- 
    ra_10037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 735_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4552_inst_ack_0, ack => zeropad3D_CP_2067_elements(735)); -- 
    -- CP-element group 736:  branch  transition  place  input  output  bypass 
    -- CP-element group 736: predecessors 
    -- CP-element group 736: 	732 
    -- CP-element group 736: successors 
    -- CP-element group 736: 	737 
    -- CP-element group 736: 	738 
    -- CP-element group 736:  members (13) 
      -- CP-element group 736: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565__exit__
      -- CP-element group 736: 	 branch_block_stmt_655/if_stmt_4566__entry__
      -- CP-element group 736: 	 branch_block_stmt_655/if_stmt_4566_else_link/$entry
      -- CP-element group 736: 	 branch_block_stmt_655/if_stmt_4566_if_link/$entry
      -- CP-element group 736: 	 branch_block_stmt_655/R_cmp1584_4567_place
      -- CP-element group 736: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/$exit
      -- CP-element group 736: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_update_completed_
      -- CP-element group 736: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_Update/$exit
      -- CP-element group 736: 	 branch_block_stmt_655/assign_stmt_4549_to_assign_stmt_4565/type_cast_4552_Update/ca
      -- CP-element group 736: 	 branch_block_stmt_655/if_stmt_4566_dead_link/$entry
      -- CP-element group 736: 	 branch_block_stmt_655/if_stmt_4566_eval_test/$entry
      -- CP-element group 736: 	 branch_block_stmt_655/if_stmt_4566_eval_test/$exit
      -- CP-element group 736: 	 branch_block_stmt_655/if_stmt_4566_eval_test/branch_req
      -- 
    ca_10042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 736_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4552_inst_ack_1, ack => zeropad3D_CP_2067_elements(736)); -- 
    branch_req_10050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(736), ack => if_stmt_4566_branch_req_0); -- 
    -- CP-element group 737:  fork  transition  place  input  output  bypass 
    -- CP-element group 737: predecessors 
    -- CP-element group 737: 	736 
    -- CP-element group 737: successors 
    -- CP-element group 737: 	753 
    -- CP-element group 737: 	754 
    -- CP-element group 737: 	756 
    -- CP-element group 737: 	758 
    -- CP-element group 737: 	760 
    -- CP-element group 737: 	762 
    -- CP-element group 737: 	764 
    -- CP-element group 737: 	766 
    -- CP-element group 737: 	768 
    -- CP-element group 737: 	771 
    -- CP-element group 737:  members (46) 
      -- CP-element group 737: 	 branch_block_stmt_655/merge_stmt_4630__exit__
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735__entry__
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_complete/req
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_update_start_
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/word_access_complete/word_0/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/word_access_complete/word_0/cr
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_update_start_
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_Update/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_complete/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_update_start_
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_update_start_
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_sample_start_
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_Update/cr
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/word_access_complete/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_Update/req
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_Update/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_Update/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_update_start_
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_update_start
      -- CP-element group 737: 	 branch_block_stmt_655/if_stmt_4566_if_link/if_choice_transition
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_Update/cr
      -- CP-element group 737: 	 branch_block_stmt_655/if_stmt_4566_if_link/$exit
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_Update/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1576_ifx_xelse1607
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_Sample/rr
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_Sample/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_Update/cr
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_update_start_
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_update_start
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_Update/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_Update/req
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_complete/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_complete/req
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_update_start_
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Update/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Update/word_access_complete/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Update/word_access_complete/word_0/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Update/word_access_complete/word_0/cr
      -- CP-element group 737: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1576_ifx_xelse1607_PhiReq/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1576_ifx_xelse1607_PhiReq/$exit
      -- CP-element group 737: 	 branch_block_stmt_655/merge_stmt_4630_PhiReqMerge
      -- CP-element group 737: 	 branch_block_stmt_655/merge_stmt_4630_PhiAck/$entry
      -- CP-element group 737: 	 branch_block_stmt_655/merge_stmt_4630_PhiAck/$exit
      -- CP-element group 737: 	 branch_block_stmt_655/merge_stmt_4630_PhiAck/dummy
      -- 
    if_choice_transition_10055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 737_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4566_branch_ack_1, ack => zeropad3D_CP_2067_elements(737)); -- 
    req_10278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => addr_of_4705_final_reg_req_1); -- 
    cr_10323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => ptr_deref_4709_load_0_req_1); -- 
    cr_10232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => type_cast_4698_inst_req_1); -- 
    req_10263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => array_obj_ref_4704_index_offset_req_1); -- 
    cr_10218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => type_cast_4634_inst_req_1); -- 
    rr_10213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => type_cast_4634_inst_req_0); -- 
    cr_10342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => type_cast_4723_inst_req_1); -- 
    req_10373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => array_obj_ref_4729_index_offset_req_1); -- 
    req_10388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => addr_of_4730_final_reg_req_1); -- 
    cr_10438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(737), ack => ptr_deref_4733_store_0_req_1); -- 
    -- CP-element group 738:  transition  place  input  bypass 
    -- CP-element group 738: predecessors 
    -- CP-element group 738: 	736 
    -- CP-element group 738: successors 
    -- CP-element group 738: 	1226 
    -- CP-element group 738:  members (5) 
      -- CP-element group 738: 	 branch_block_stmt_655/if_stmt_4566_else_link/else_choice_transition
      -- CP-element group 738: 	 branch_block_stmt_655/if_stmt_4566_else_link/$exit
      -- CP-element group 738: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1576_ifx_xthen1586
      -- CP-element group 738: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1576_ifx_xthen1586_PhiReq/$entry
      -- CP-element group 738: 	 branch_block_stmt_655/lorx_xlhsx_xfalse1576_ifx_xthen1586_PhiReq/$exit
      -- 
    else_choice_transition_10059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 738_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4566_branch_ack_0, ack => zeropad3D_CP_2067_elements(738)); -- 
    -- CP-element group 739:  transition  input  bypass 
    -- CP-element group 739: predecessors 
    -- CP-element group 739: 	1226 
    -- CP-element group 739: successors 
    -- CP-element group 739:  members (3) 
      -- CP-element group 739: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_Sample/ra
      -- CP-element group 739: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_Sample/$exit
      -- CP-element group 739: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_sample_completed_
      -- 
    ra_10073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 739_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4576_inst_ack_0, ack => zeropad3D_CP_2067_elements(739)); -- 
    -- CP-element group 740:  transition  input  bypass 
    -- CP-element group 740: predecessors 
    -- CP-element group 740: 	1226 
    -- CP-element group 740: successors 
    -- CP-element group 740: 	743 
    -- CP-element group 740:  members (3) 
      -- CP-element group 740: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_Update/ca
      -- CP-element group 740: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_Update/$exit
      -- CP-element group 740: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_update_completed_
      -- 
    ca_10078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 740_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4576_inst_ack_1, ack => zeropad3D_CP_2067_elements(740)); -- 
    -- CP-element group 741:  transition  input  bypass 
    -- CP-element group 741: predecessors 
    -- CP-element group 741: 	1226 
    -- CP-element group 741: successors 
    -- CP-element group 741:  members (3) 
      -- CP-element group 741: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_Sample/ra
      -- CP-element group 741: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_Sample/$exit
      -- CP-element group 741: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_sample_completed_
      -- 
    ra_10087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 741_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4581_inst_ack_0, ack => zeropad3D_CP_2067_elements(741)); -- 
    -- CP-element group 742:  transition  input  bypass 
    -- CP-element group 742: predecessors 
    -- CP-element group 742: 	1226 
    -- CP-element group 742: successors 
    -- CP-element group 742: 	743 
    -- CP-element group 742:  members (3) 
      -- CP-element group 742: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_Update/ca
      -- CP-element group 742: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_Update/$exit
      -- CP-element group 742: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_update_completed_
      -- 
    ca_10092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 742_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4581_inst_ack_1, ack => zeropad3D_CP_2067_elements(742)); -- 
    -- CP-element group 743:  join  transition  output  bypass 
    -- CP-element group 743: predecessors 
    -- CP-element group 743: 	740 
    -- CP-element group 743: 	742 
    -- CP-element group 743: successors 
    -- CP-element group 743: 	744 
    -- CP-element group 743:  members (3) 
      -- CP-element group 743: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_sample_start_
      -- CP-element group 743: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_Sample/rr
      -- CP-element group 743: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_Sample/$entry
      -- 
    rr_10100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(743), ack => type_cast_4615_inst_req_0); -- 
    zeropad3D_cp_element_group_743: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_743"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(740) & zeropad3D_CP_2067_elements(742);
      gj_zeropad3D_cp_element_group_743 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(743), clk => clk, reset => reset); --
    end block;
    -- CP-element group 744:  transition  input  bypass 
    -- CP-element group 744: predecessors 
    -- CP-element group 744: 	743 
    -- CP-element group 744: successors 
    -- CP-element group 744:  members (3) 
      -- CP-element group 744: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_sample_completed_
      -- CP-element group 744: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_Sample/ra
      -- CP-element group 744: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_Sample/$exit
      -- 
    ra_10101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 744_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4615_inst_ack_0, ack => zeropad3D_CP_2067_elements(744)); -- 
    -- CP-element group 745:  transition  input  output  bypass 
    -- CP-element group 745: predecessors 
    -- CP-element group 745: 	1226 
    -- CP-element group 745: successors 
    -- CP-element group 745: 	746 
    -- CP-element group 745:  members (16) 
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_resized_1
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_scaled_1
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_scale_1/scale_rename_req
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_scale_1/$exit
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_scale_1/$entry
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_resize_1/index_resize_ack
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_resize_1/index_resize_req
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_resize_1/$exit
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_Update/ca
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_resize_1/$entry
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_computed_1
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_Update/$exit
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_Sample/req
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_update_completed_
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_Sample/$entry
      -- CP-element group 745: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_index_scale_1/scale_rename_ack
      -- 
    ca_10106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 745_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4615_inst_ack_1, ack => zeropad3D_CP_2067_elements(745)); -- 
    req_10131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(745), ack => array_obj_ref_4621_index_offset_req_0); -- 
    -- CP-element group 746:  transition  input  bypass 
    -- CP-element group 746: predecessors 
    -- CP-element group 746: 	745 
    -- CP-element group 746: successors 
    -- CP-element group 746: 	752 
    -- CP-element group 746:  members (3) 
      -- CP-element group 746: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_Sample/ack
      -- CP-element group 746: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_Sample/$exit
      -- CP-element group 746: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_sample_complete
      -- 
    ack_10132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 746_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4621_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(746)); -- 
    -- CP-element group 747:  transition  input  output  bypass 
    -- CP-element group 747: predecessors 
    -- CP-element group 747: 	1226 
    -- CP-element group 747: successors 
    -- CP-element group 747: 	748 
    -- CP-element group 747:  members (11) 
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_offset_calculated
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_root_address_calculated
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_sample_start_
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_request/req
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_request/$entry
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_base_plus_offset/sum_rename_ack
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_base_plus_offset/sum_rename_req
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_base_plus_offset/$exit
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_base_plus_offset/$entry
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_Update/ack
      -- CP-element group 747: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_Update/$exit
      -- 
    ack_10137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 747_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4621_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(747)); -- 
    req_10146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(747), ack => addr_of_4622_final_reg_req_0); -- 
    -- CP-element group 748:  transition  input  bypass 
    -- CP-element group 748: predecessors 
    -- CP-element group 748: 	747 
    -- CP-element group 748: successors 
    -- CP-element group 748:  members (3) 
      -- CP-element group 748: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_sample_completed_
      -- CP-element group 748: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_request/ack
      -- CP-element group 748: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_request/$exit
      -- 
    ack_10147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 748_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4622_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(748)); -- 
    -- CP-element group 749:  join  fork  transition  input  output  bypass 
    -- CP-element group 749: predecessors 
    -- CP-element group 749: 	1226 
    -- CP-element group 749: successors 
    -- CP-element group 749: 	750 
    -- CP-element group 749:  members (28) 
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/word_access_start/word_0/$entry
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/word_access_start/word_0/rr
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/word_access_start/$entry
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/ptr_deref_4625_Split/split_ack
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/ptr_deref_4625_Split/split_req
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/ptr_deref_4625_Split/$exit
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/ptr_deref_4625_Split/$entry
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/$entry
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_word_addrgen/root_register_ack
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_word_addrgen/root_register_req
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_word_addrgen/$exit
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_word_addrgen/$entry
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_plus_offset/sum_rename_ack
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_plus_offset/sum_rename_req
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_plus_offset/$exit
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_plus_offset/$entry
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_addr_resize/base_resize_ack
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_addr_resize/base_resize_req
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_addr_resize/$exit
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_addr_resize/$entry
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_address_resized
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_root_address_calculated
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_word_address_calculated
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_update_completed_
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_base_address_calculated
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_sample_start_
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_complete/ack
      -- CP-element group 749: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_complete/$exit
      -- 
    ack_10152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 749_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4622_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(749)); -- 
    rr_10190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(749), ack => ptr_deref_4625_store_0_req_0); -- 
    -- CP-element group 750:  transition  input  bypass 
    -- CP-element group 750: predecessors 
    -- CP-element group 750: 	749 
    -- CP-element group 750: successors 
    -- CP-element group 750:  members (5) 
      -- CP-element group 750: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/word_access_start/word_0/$exit
      -- CP-element group 750: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/word_access_start/word_0/ra
      -- CP-element group 750: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/word_access_start/$exit
      -- CP-element group 750: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Sample/$exit
      -- CP-element group 750: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_sample_completed_
      -- 
    ra_10191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 750_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4625_store_0_ack_0, ack => zeropad3D_CP_2067_elements(750)); -- 
    -- CP-element group 751:  transition  input  bypass 
    -- CP-element group 751: predecessors 
    -- CP-element group 751: 	1226 
    -- CP-element group 751: successors 
    -- CP-element group 751: 	752 
    -- CP-element group 751:  members (5) 
      -- CP-element group 751: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Update/word_access_complete/word_0/ca
      -- CP-element group 751: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_update_completed_
      -- CP-element group 751: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Update/word_access_complete/word_0/$exit
      -- CP-element group 751: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Update/word_access_complete/$exit
      -- CP-element group 751: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Update/$exit
      -- 
    ca_10202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 751_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4625_store_0_ack_1, ack => zeropad3D_CP_2067_elements(751)); -- 
    -- CP-element group 752:  join  transition  place  bypass 
    -- CP-element group 752: predecessors 
    -- CP-element group 752: 	746 
    -- CP-element group 752: 	751 
    -- CP-element group 752: successors 
    -- CP-element group 752: 	1227 
    -- CP-element group 752:  members (5) 
      -- CP-element group 752: 	 branch_block_stmt_655/ifx_xthen1586_ifx_xend1655
      -- CP-element group 752: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628__exit__
      -- CP-element group 752: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/$exit
      -- CP-element group 752: 	 branch_block_stmt_655/ifx_xthen1586_ifx_xend1655_PhiReq/$entry
      -- CP-element group 752: 	 branch_block_stmt_655/ifx_xthen1586_ifx_xend1655_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_752: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_752"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(746) & zeropad3D_CP_2067_elements(751);
      gj_zeropad3D_cp_element_group_752 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(752), clk => clk, reset => reset); --
    end block;
    -- CP-element group 753:  transition  input  bypass 
    -- CP-element group 753: predecessors 
    -- CP-element group 753: 	737 
    -- CP-element group 753: successors 
    -- CP-element group 753:  members (3) 
      -- CP-element group 753: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_sample_completed_
      -- CP-element group 753: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_Sample/ra
      -- CP-element group 753: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_Sample/$exit
      -- 
    ra_10214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 753_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4634_inst_ack_0, ack => zeropad3D_CP_2067_elements(753)); -- 
    -- CP-element group 754:  fork  transition  input  output  bypass 
    -- CP-element group 754: predecessors 
    -- CP-element group 754: 	737 
    -- CP-element group 754: successors 
    -- CP-element group 754: 	755 
    -- CP-element group 754: 	763 
    -- CP-element group 754:  members (9) 
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_update_completed_
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_Sample/rr
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_sample_start_
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_Sample/$entry
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_Sample/rr
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_Sample/$entry
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_sample_start_
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_Update/ca
      -- CP-element group 754: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4634_Update/$exit
      -- 
    ca_10219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 754_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4634_inst_ack_1, ack => zeropad3D_CP_2067_elements(754)); -- 
    rr_10227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(754), ack => type_cast_4698_inst_req_0); -- 
    rr_10337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(754), ack => type_cast_4723_inst_req_0); -- 
    -- CP-element group 755:  transition  input  bypass 
    -- CP-element group 755: predecessors 
    -- CP-element group 755: 	754 
    -- CP-element group 755: successors 
    -- CP-element group 755:  members (3) 
      -- CP-element group 755: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_Sample/ra
      -- CP-element group 755: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_Sample/$exit
      -- CP-element group 755: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_sample_completed_
      -- 
    ra_10228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 755_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4698_inst_ack_0, ack => zeropad3D_CP_2067_elements(755)); -- 
    -- CP-element group 756:  transition  input  output  bypass 
    -- CP-element group 756: predecessors 
    -- CP-element group 756: 	737 
    -- CP-element group 756: successors 
    -- CP-element group 756: 	757 
    -- CP-element group 756:  members (16) 
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_resize_1/index_resize_ack
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_resize_1/index_resize_req
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_resize_1/$exit
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_resize_1/$entry
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_computed_1
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_scaled_1
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_resized_1
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_Update/ca
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_Update/$exit
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4698_update_completed_
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_Sample/req
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_Sample/$entry
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_scale_1/scale_rename_ack
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_scale_1/scale_rename_req
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_scale_1/$exit
      -- CP-element group 756: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_index_scale_1/$entry
      -- 
    ca_10233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 756_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4698_inst_ack_1, ack => zeropad3D_CP_2067_elements(756)); -- 
    req_10258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(756), ack => array_obj_ref_4704_index_offset_req_0); -- 
    -- CP-element group 757:  transition  input  bypass 
    -- CP-element group 757: predecessors 
    -- CP-element group 757: 	756 
    -- CP-element group 757: successors 
    -- CP-element group 757: 	772 
    -- CP-element group 757:  members (3) 
      -- CP-element group 757: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_Sample/ack
      -- CP-element group 757: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_Sample/$exit
      -- CP-element group 757: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_sample_complete
      -- 
    ack_10259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 757_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4704_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(757)); -- 
    -- CP-element group 758:  transition  input  output  bypass 
    -- CP-element group 758: predecessors 
    -- CP-element group 758: 	737 
    -- CP-element group 758: successors 
    -- CP-element group 758: 	759 
    -- CP-element group 758:  members (11) 
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_request/req
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_request/$entry
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_base_plus_offset/sum_rename_ack
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_base_plus_offset/sum_rename_req
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_base_plus_offset/$exit
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_offset_calculated
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_root_address_calculated
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_base_plus_offset/$entry
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_sample_start_
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_Update/ack
      -- CP-element group 758: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4704_final_index_sum_regn_Update/$exit
      -- 
    ack_10264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 758_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4704_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(758)); -- 
    req_10273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(758), ack => addr_of_4705_final_reg_req_0); -- 
    -- CP-element group 759:  transition  input  bypass 
    -- CP-element group 759: predecessors 
    -- CP-element group 759: 	758 
    -- CP-element group 759: successors 
    -- CP-element group 759:  members (3) 
      -- CP-element group 759: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_request/ack
      -- CP-element group 759: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_request/$exit
      -- CP-element group 759: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_sample_completed_
      -- 
    ack_10274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 759_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4705_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(759)); -- 
    -- CP-element group 760:  join  fork  transition  input  output  bypass 
    -- CP-element group 760: predecessors 
    -- CP-element group 760: 	737 
    -- CP-element group 760: successors 
    -- CP-element group 760: 	761 
    -- CP-element group 760:  members (24) 
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_complete/ack
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_sample_start_
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_complete/$exit
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_address_resized
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Sample/word_access_start/word_0/$entry
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_root_address_calculated
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4705_update_completed_
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_word_address_calculated
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Sample/word_access_start/$entry
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Sample/word_access_start/word_0/rr
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_address_calculated
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Sample/$entry
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_word_addrgen/root_register_ack
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_word_addrgen/root_register_req
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_word_addrgen/$exit
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_word_addrgen/$entry
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_plus_offset/sum_rename_ack
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_plus_offset/sum_rename_req
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_plus_offset/$exit
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_plus_offset/$entry
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_addr_resize/base_resize_ack
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_addr_resize/base_resize_req
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_addr_resize/$exit
      -- CP-element group 760: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_base_addr_resize/$entry
      -- 
    ack_10279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 760_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4705_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(760)); -- 
    rr_10312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(760), ack => ptr_deref_4709_load_0_req_0); -- 
    -- CP-element group 761:  transition  input  bypass 
    -- CP-element group 761: predecessors 
    -- CP-element group 761: 	760 
    -- CP-element group 761: successors 
    -- CP-element group 761:  members (5) 
      -- CP-element group 761: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_sample_completed_
      -- CP-element group 761: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Sample/word_access_start/word_0/ra
      -- CP-element group 761: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Sample/word_access_start/word_0/$exit
      -- CP-element group 761: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Sample/word_access_start/$exit
      -- CP-element group 761: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Sample/$exit
      -- 
    ra_10313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 761_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4709_load_0_ack_0, ack => zeropad3D_CP_2067_elements(761)); -- 
    -- CP-element group 762:  transition  input  bypass 
    -- CP-element group 762: predecessors 
    -- CP-element group 762: 	737 
    -- CP-element group 762: successors 
    -- CP-element group 762: 	769 
    -- CP-element group 762:  members (9) 
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/word_access_complete/word_0/$exit
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/word_access_complete/$exit
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/$exit
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/ptr_deref_4709_Merge/merge_ack
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/ptr_deref_4709_Merge/merge_req
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/ptr_deref_4709_Merge/$exit
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/ptr_deref_4709_Merge/$entry
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_Update/word_access_complete/word_0/ca
      -- CP-element group 762: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4709_update_completed_
      -- 
    ca_10324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 762_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4709_load_0_ack_1, ack => zeropad3D_CP_2067_elements(762)); -- 
    -- CP-element group 763:  transition  input  bypass 
    -- CP-element group 763: predecessors 
    -- CP-element group 763: 	754 
    -- CP-element group 763: successors 
    -- CP-element group 763:  members (3) 
      -- CP-element group 763: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_Sample/ra
      -- CP-element group 763: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_sample_completed_
      -- CP-element group 763: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_Sample/$exit
      -- 
    ra_10338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 763_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4723_inst_ack_0, ack => zeropad3D_CP_2067_elements(763)); -- 
    -- CP-element group 764:  transition  input  output  bypass 
    -- CP-element group 764: predecessors 
    -- CP-element group 764: 	737 
    -- CP-element group 764: successors 
    -- CP-element group 764: 	765 
    -- CP-element group 764:  members (16) 
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_Update/$exit
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_update_completed_
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/type_cast_4723_Update/ca
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_resized_1
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_scaled_1
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_computed_1
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_resize_1/$entry
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_resize_1/$exit
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_resize_1/index_resize_req
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_resize_1/index_resize_ack
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_scale_1/$entry
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_scale_1/$exit
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_scale_1/scale_rename_req
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_index_scale_1/scale_rename_ack
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_Sample/$entry
      -- CP-element group 764: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_Sample/req
      -- 
    ca_10343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 764_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4723_inst_ack_1, ack => zeropad3D_CP_2067_elements(764)); -- 
    req_10368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(764), ack => array_obj_ref_4729_index_offset_req_0); -- 
    -- CP-element group 765:  transition  input  bypass 
    -- CP-element group 765: predecessors 
    -- CP-element group 765: 	764 
    -- CP-element group 765: successors 
    -- CP-element group 765: 	772 
    -- CP-element group 765:  members (3) 
      -- CP-element group 765: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_sample_complete
      -- CP-element group 765: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_Sample/$exit
      -- CP-element group 765: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_Sample/ack
      -- 
    ack_10369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 765_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4729_index_offset_ack_0, ack => zeropad3D_CP_2067_elements(765)); -- 
    -- CP-element group 766:  transition  input  output  bypass 
    -- CP-element group 766: predecessors 
    -- CP-element group 766: 	737 
    -- CP-element group 766: successors 
    -- CP-element group 766: 	767 
    -- CP-element group 766:  members (11) 
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_request/$entry
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_sample_start_
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_root_address_calculated
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_offset_calculated
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_Update/$exit
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_final_index_sum_regn_Update/ack
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_base_plus_offset/$entry
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_base_plus_offset/$exit
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_base_plus_offset/sum_rename_req
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/array_obj_ref_4729_base_plus_offset/sum_rename_ack
      -- CP-element group 766: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_request/req
      -- 
    ack_10374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 766_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4729_index_offset_ack_1, ack => zeropad3D_CP_2067_elements(766)); -- 
    req_10383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(766), ack => addr_of_4730_final_reg_req_0); -- 
    -- CP-element group 767:  transition  input  bypass 
    -- CP-element group 767: predecessors 
    -- CP-element group 767: 	766 
    -- CP-element group 767: successors 
    -- CP-element group 767:  members (3) 
      -- CP-element group 767: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_sample_completed_
      -- CP-element group 767: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_request/$exit
      -- CP-element group 767: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_request/ack
      -- 
    ack_10384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 767_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4730_final_reg_ack_0, ack => zeropad3D_CP_2067_elements(767)); -- 
    -- CP-element group 768:  fork  transition  input  bypass 
    -- CP-element group 768: predecessors 
    -- CP-element group 768: 	737 
    -- CP-element group 768: successors 
    -- CP-element group 768: 	769 
    -- CP-element group 768:  members (19) 
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_update_completed_
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_complete/$exit
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/addr_of_4730_complete/ack
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_address_calculated
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_word_address_calculated
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_root_address_calculated
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_address_resized
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_addr_resize/$entry
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_addr_resize/$exit
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_addr_resize/base_resize_req
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_addr_resize/base_resize_ack
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_plus_offset/$entry
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_plus_offset/$exit
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_plus_offset/sum_rename_req
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_base_plus_offset/sum_rename_ack
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_word_addrgen/$entry
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_word_addrgen/$exit
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_word_addrgen/root_register_req
      -- CP-element group 768: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_word_addrgen/root_register_ack
      -- 
    ack_10389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 768_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4730_final_reg_ack_1, ack => zeropad3D_CP_2067_elements(768)); -- 
    -- CP-element group 769:  join  transition  output  bypass 
    -- CP-element group 769: predecessors 
    -- CP-element group 769: 	762 
    -- CP-element group 769: 	768 
    -- CP-element group 769: successors 
    -- CP-element group 769: 	770 
    -- CP-element group 769:  members (9) 
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_sample_start_
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/$entry
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/ptr_deref_4733_Split/$entry
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/ptr_deref_4733_Split/$exit
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/ptr_deref_4733_Split/split_req
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/ptr_deref_4733_Split/split_ack
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/word_access_start/$entry
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/word_access_start/word_0/$entry
      -- CP-element group 769: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/word_access_start/word_0/rr
      -- 
    rr_10427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(769), ack => ptr_deref_4733_store_0_req_0); -- 
    zeropad3D_cp_element_group_769: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_769"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(762) & zeropad3D_CP_2067_elements(768);
      gj_zeropad3D_cp_element_group_769 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(769), clk => clk, reset => reset); --
    end block;
    -- CP-element group 770:  transition  input  bypass 
    -- CP-element group 770: predecessors 
    -- CP-element group 770: 	769 
    -- CP-element group 770: successors 
    -- CP-element group 770:  members (5) 
      -- CP-element group 770: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_sample_completed_
      -- CP-element group 770: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/$exit
      -- CP-element group 770: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/word_access_start/$exit
      -- CP-element group 770: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/word_access_start/word_0/$exit
      -- CP-element group 770: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Sample/word_access_start/word_0/ra
      -- 
    ra_10428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 770_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4733_store_0_ack_0, ack => zeropad3D_CP_2067_elements(770)); -- 
    -- CP-element group 771:  transition  input  bypass 
    -- CP-element group 771: predecessors 
    -- CP-element group 771: 	737 
    -- CP-element group 771: successors 
    -- CP-element group 771: 	772 
    -- CP-element group 771:  members (5) 
      -- CP-element group 771: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_update_completed_
      -- CP-element group 771: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Update/$exit
      -- CP-element group 771: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Update/word_access_complete/$exit
      -- CP-element group 771: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Update/word_access_complete/word_0/$exit
      -- CP-element group 771: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/ptr_deref_4733_Update/word_access_complete/word_0/ca
      -- 
    ca_10439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 771_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4733_store_0_ack_1, ack => zeropad3D_CP_2067_elements(771)); -- 
    -- CP-element group 772:  join  transition  place  bypass 
    -- CP-element group 772: predecessors 
    -- CP-element group 772: 	757 
    -- CP-element group 772: 	765 
    -- CP-element group 772: 	771 
    -- CP-element group 772: successors 
    -- CP-element group 772: 	1227 
    -- CP-element group 772:  members (5) 
      -- CP-element group 772: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735__exit__
      -- CP-element group 772: 	 branch_block_stmt_655/ifx_xelse1607_ifx_xend1655
      -- CP-element group 772: 	 branch_block_stmt_655/assign_stmt_4635_to_assign_stmt_4735/$exit
      -- CP-element group 772: 	 branch_block_stmt_655/ifx_xelse1607_ifx_xend1655_PhiReq/$entry
      -- CP-element group 772: 	 branch_block_stmt_655/ifx_xelse1607_ifx_xend1655_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_772: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_772"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(757) & zeropad3D_CP_2067_elements(765) & zeropad3D_CP_2067_elements(771);
      gj_zeropad3D_cp_element_group_772 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(772), clk => clk, reset => reset); --
    end block;
    -- CP-element group 773:  transition  input  bypass 
    -- CP-element group 773: predecessors 
    -- CP-element group 773: 	1227 
    -- CP-element group 773: successors 
    -- CP-element group 773:  members (3) 
      -- CP-element group 773: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_sample_completed_
      -- CP-element group 773: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_Sample/$exit
      -- CP-element group 773: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_Sample/ra
      -- 
    ra_10451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 773_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4741_inst_ack_0, ack => zeropad3D_CP_2067_elements(773)); -- 
    -- CP-element group 774:  branch  transition  place  input  output  bypass 
    -- CP-element group 774: predecessors 
    -- CP-element group 774: 	1227 
    -- CP-element group 774: successors 
    -- CP-element group 774: 	775 
    -- CP-element group 774: 	776 
    -- CP-element group 774:  members (13) 
      -- CP-element group 774: 	 branch_block_stmt_655/if_stmt_4756__entry__
      -- CP-element group 774: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755__exit__
      -- CP-element group 774: 	 branch_block_stmt_655/R_cmp1663_4757_place
      -- CP-element group 774: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/$exit
      -- CP-element group 774: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_update_completed_
      -- CP-element group 774: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_Update/$exit
      -- CP-element group 774: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_Update/ca
      -- CP-element group 774: 	 branch_block_stmt_655/if_stmt_4756_dead_link/$entry
      -- CP-element group 774: 	 branch_block_stmt_655/if_stmt_4756_eval_test/$entry
      -- CP-element group 774: 	 branch_block_stmt_655/if_stmt_4756_eval_test/$exit
      -- CP-element group 774: 	 branch_block_stmt_655/if_stmt_4756_eval_test/branch_req
      -- CP-element group 774: 	 branch_block_stmt_655/if_stmt_4756_if_link/$entry
      -- CP-element group 774: 	 branch_block_stmt_655/if_stmt_4756_else_link/$entry
      -- 
    ca_10456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 774_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4741_inst_ack_1, ack => zeropad3D_CP_2067_elements(774)); -- 
    branch_req_10464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(774), ack => if_stmt_4756_branch_req_0); -- 
    -- CP-element group 775:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 775: predecessors 
    -- CP-element group 775: 	774 
    -- CP-element group 775: successors 
    -- CP-element group 775: 	1236 
    -- CP-element group 775: 	1237 
    -- CP-element group 775: 	1239 
    -- CP-element group 775: 	1240 
    -- CP-element group 775: 	1242 
    -- CP-element group 775: 	1243 
    -- CP-element group 775:  members (40) 
      -- CP-element group 775: 	 branch_block_stmt_655/assign_stmt_4768__exit__
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705
      -- CP-element group 775: 	 branch_block_stmt_655/merge_stmt_4762__exit__
      -- CP-element group 775: 	 branch_block_stmt_655/assign_stmt_4768__entry__
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xend1655_ifx_xthen1665
      -- CP-element group 775: 	 branch_block_stmt_655/if_stmt_4756_if_link/$exit
      -- CP-element group 775: 	 branch_block_stmt_655/if_stmt_4756_if_link/if_choice_transition
      -- CP-element group 775: 	 branch_block_stmt_655/assign_stmt_4768/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/assign_stmt_4768/$exit
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xend1655_ifx_xthen1665_PhiReq/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xend1655_ifx_xthen1665_PhiReq/$exit
      -- CP-element group 775: 	 branch_block_stmt_655/merge_stmt_4762_PhiReqMerge
      -- CP-element group 775: 	 branch_block_stmt_655/merge_stmt_4762_PhiAck/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/merge_stmt_4762_PhiAck/$exit
      -- CP-element group 775: 	 branch_block_stmt_655/merge_stmt_4762_PhiAck/dummy
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/Sample/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/Sample/rr
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/Update/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/Update/cr
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/Sample/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/Sample/rr
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/Update/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/Update/cr
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/Sample/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/Sample/rr
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/Update/$entry
      -- CP-element group 775: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/Update/cr
      -- 
    if_choice_transition_10469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 775_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4756_branch_ack_1, ack => zeropad3D_CP_2067_elements(775)); -- 
    rr_13936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(775), ack => type_cast_4859_inst_req_0); -- 
    cr_13941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(775), ack => type_cast_4859_inst_req_1); -- 
    rr_13959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(775), ack => type_cast_4849_inst_req_0); -- 
    cr_13964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(775), ack => type_cast_4849_inst_req_1); -- 
    rr_13982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(775), ack => type_cast_4853_inst_req_0); -- 
    cr_13987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(775), ack => type_cast_4853_inst_req_1); -- 
    -- CP-element group 776:  fork  transition  place  input  output  bypass 
    -- CP-element group 776: predecessors 
    -- CP-element group 776: 	774 
    -- CP-element group 776: successors 
    -- CP-element group 776: 	777 
    -- CP-element group 776: 	778 
    -- CP-element group 776: 	779 
    -- CP-element group 776: 	780 
    -- CP-element group 776: 	782 
    -- CP-element group 776: 	785 
    -- CP-element group 776: 	787 
    -- CP-element group 776: 	788 
    -- CP-element group 776: 	789 
    -- CP-element group 776: 	791 
    -- CP-element group 776:  members (54) 
      -- CP-element group 776: 	 branch_block_stmt_655/merge_stmt_4770__exit__
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835__entry__
      -- CP-element group 776: 	 branch_block_stmt_655/ifx_xend1655_ifx_xelse1670
      -- CP-element group 776: 	 branch_block_stmt_655/if_stmt_4756_else_link/$exit
      -- CP-element group 776: 	 branch_block_stmt_655/if_stmt_4756_else_link/else_choice_transition
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_sample_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_update_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_Sample/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_Sample/rr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_Update/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_Update/cr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_sample_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_update_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_word_address_calculated
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_root_address_calculated
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Sample/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Sample/word_access_start/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Sample/word_access_start/word_0/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Sample/word_access_start/word_0/rr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/word_access_complete/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/word_access_complete/word_0/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/word_access_complete/word_0/cr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_update_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_Update/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_Update/cr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_update_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_Update/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_Update/cr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_update_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_Update/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_Update/cr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_sample_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_update_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_word_address_calculated
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_root_address_calculated
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Sample/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Sample/word_access_start/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Sample/word_access_start/word_0/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Sample/word_access_start/word_0/rr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/word_access_complete/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/word_access_complete/word_0/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/word_access_complete/word_0/cr
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_update_start_
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_Update/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_Update/cr
      -- CP-element group 776: 	 branch_block_stmt_655/ifx_xend1655_ifx_xelse1670_PhiReq/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/ifx_xend1655_ifx_xelse1670_PhiReq/$exit
      -- CP-element group 776: 	 branch_block_stmt_655/merge_stmt_4770_PhiReqMerge
      -- CP-element group 776: 	 branch_block_stmt_655/merge_stmt_4770_PhiAck/$entry
      -- CP-element group 776: 	 branch_block_stmt_655/merge_stmt_4770_PhiAck/$exit
      -- CP-element group 776: 	 branch_block_stmt_655/merge_stmt_4770_PhiAck/dummy
      -- 
    else_choice_transition_10473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 776_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4756_branch_ack_0, ack => zeropad3D_CP_2067_elements(776)); -- 
    rr_10489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => type_cast_4780_inst_req_0); -- 
    cr_10494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => type_cast_4780_inst_req_1); -- 
    rr_10511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => LOAD_col_high_4783_load_0_req_0); -- 
    cr_10522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => LOAD_col_high_4783_load_0_req_1); -- 
    cr_10541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => type_cast_4787_inst_req_1); -- 
    cr_10555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => type_cast_4801_inst_req_1); -- 
    cr_10569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => type_cast_4817_inst_req_1); -- 
    rr_10586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => LOAD_row_high_4820_load_0_req_0); -- 
    cr_10597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => LOAD_row_high_4820_load_0_req_1); -- 
    cr_10616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(776), ack => type_cast_4824_inst_req_1); -- 
    -- CP-element group 777:  transition  input  bypass 
    -- CP-element group 777: predecessors 
    -- CP-element group 777: 	776 
    -- CP-element group 777: successors 
    -- CP-element group 777:  members (3) 
      -- CP-element group 777: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_sample_completed_
      -- CP-element group 777: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_Sample/$exit
      -- CP-element group 777: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_Sample/ra
      -- 
    ra_10490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 777_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4780_inst_ack_0, ack => zeropad3D_CP_2067_elements(777)); -- 
    -- CP-element group 778:  transition  input  bypass 
    -- CP-element group 778: predecessors 
    -- CP-element group 778: 	776 
    -- CP-element group 778: successors 
    -- CP-element group 778: 	783 
    -- CP-element group 778:  members (3) 
      -- CP-element group 778: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_update_completed_
      -- CP-element group 778: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_Update/$exit
      -- CP-element group 778: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4780_Update/ca
      -- 
    ca_10495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 778_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4780_inst_ack_1, ack => zeropad3D_CP_2067_elements(778)); -- 
    -- CP-element group 779:  transition  input  bypass 
    -- CP-element group 779: predecessors 
    -- CP-element group 779: 	776 
    -- CP-element group 779: successors 
    -- CP-element group 779:  members (5) 
      -- CP-element group 779: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_sample_completed_
      -- CP-element group 779: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Sample/$exit
      -- CP-element group 779: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Sample/word_access_start/$exit
      -- CP-element group 779: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Sample/word_access_start/word_0/$exit
      -- CP-element group 779: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Sample/word_access_start/word_0/ra
      -- 
    ra_10512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 779_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4783_load_0_ack_0, ack => zeropad3D_CP_2067_elements(779)); -- 
    -- CP-element group 780:  transition  input  output  bypass 
    -- CP-element group 780: predecessors 
    -- CP-element group 780: 	776 
    -- CP-element group 780: successors 
    -- CP-element group 780: 	781 
    -- CP-element group 780:  members (12) 
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_update_completed_
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/$exit
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/word_access_complete/$exit
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/word_access_complete/word_0/$exit
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/word_access_complete/word_0/ca
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/LOAD_col_high_4783_Merge/$entry
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/LOAD_col_high_4783_Merge/$exit
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/LOAD_col_high_4783_Merge/merge_req
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_col_high_4783_Update/LOAD_col_high_4783_Merge/merge_ack
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_sample_start_
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_Sample/$entry
      -- CP-element group 780: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_Sample/rr
      -- 
    ca_10523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 780_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4783_load_0_ack_1, ack => zeropad3D_CP_2067_elements(780)); -- 
    rr_10536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(780), ack => type_cast_4787_inst_req_0); -- 
    -- CP-element group 781:  transition  input  bypass 
    -- CP-element group 781: predecessors 
    -- CP-element group 781: 	780 
    -- CP-element group 781: successors 
    -- CP-element group 781:  members (3) 
      -- CP-element group 781: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_sample_completed_
      -- CP-element group 781: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_Sample/$exit
      -- CP-element group 781: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_Sample/ra
      -- 
    ra_10537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 781_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4787_inst_ack_0, ack => zeropad3D_CP_2067_elements(781)); -- 
    -- CP-element group 782:  transition  input  bypass 
    -- CP-element group 782: predecessors 
    -- CP-element group 782: 	776 
    -- CP-element group 782: successors 
    -- CP-element group 782: 	783 
    -- CP-element group 782:  members (3) 
      -- CP-element group 782: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_update_completed_
      -- CP-element group 782: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_Update/$exit
      -- CP-element group 782: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4787_Update/ca
      -- 
    ca_10542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 782_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4787_inst_ack_1, ack => zeropad3D_CP_2067_elements(782)); -- 
    -- CP-element group 783:  join  transition  output  bypass 
    -- CP-element group 783: predecessors 
    -- CP-element group 783: 	778 
    -- CP-element group 783: 	782 
    -- CP-element group 783: successors 
    -- CP-element group 783: 	784 
    -- CP-element group 783:  members (3) 
      -- CP-element group 783: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_sample_start_
      -- CP-element group 783: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_Sample/$entry
      -- CP-element group 783: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_Sample/rr
      -- 
    rr_10550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(783), ack => type_cast_4801_inst_req_0); -- 
    zeropad3D_cp_element_group_783: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_783"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(778) & zeropad3D_CP_2067_elements(782);
      gj_zeropad3D_cp_element_group_783 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(783), clk => clk, reset => reset); --
    end block;
    -- CP-element group 784:  transition  input  bypass 
    -- CP-element group 784: predecessors 
    -- CP-element group 784: 	783 
    -- CP-element group 784: successors 
    -- CP-element group 784:  members (3) 
      -- CP-element group 784: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_sample_completed_
      -- CP-element group 784: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_Sample/$exit
      -- CP-element group 784: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_Sample/ra
      -- 
    ra_10551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 784_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4801_inst_ack_0, ack => zeropad3D_CP_2067_elements(784)); -- 
    -- CP-element group 785:  transition  input  output  bypass 
    -- CP-element group 785: predecessors 
    -- CP-element group 785: 	776 
    -- CP-element group 785: successors 
    -- CP-element group 785: 	786 
    -- CP-element group 785:  members (6) 
      -- CP-element group 785: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_update_completed_
      -- CP-element group 785: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_Update/$exit
      -- CP-element group 785: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4801_Update/ca
      -- CP-element group 785: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_sample_start_
      -- CP-element group 785: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_Sample/$entry
      -- CP-element group 785: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_Sample/rr
      -- 
    ca_10556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 785_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4801_inst_ack_1, ack => zeropad3D_CP_2067_elements(785)); -- 
    rr_10564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(785), ack => type_cast_4817_inst_req_0); -- 
    -- CP-element group 786:  transition  input  bypass 
    -- CP-element group 786: predecessors 
    -- CP-element group 786: 	785 
    -- CP-element group 786: successors 
    -- CP-element group 786:  members (3) 
      -- CP-element group 786: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_sample_completed_
      -- CP-element group 786: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_Sample/$exit
      -- CP-element group 786: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_Sample/ra
      -- 
    ra_10565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 786_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4817_inst_ack_0, ack => zeropad3D_CP_2067_elements(786)); -- 
    -- CP-element group 787:  transition  input  bypass 
    -- CP-element group 787: predecessors 
    -- CP-element group 787: 	776 
    -- CP-element group 787: successors 
    -- CP-element group 787: 	792 
    -- CP-element group 787:  members (3) 
      -- CP-element group 787: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_update_completed_
      -- CP-element group 787: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_Update/$exit
      -- CP-element group 787: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4817_Update/ca
      -- 
    ca_10570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 787_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4817_inst_ack_1, ack => zeropad3D_CP_2067_elements(787)); -- 
    -- CP-element group 788:  transition  input  bypass 
    -- CP-element group 788: predecessors 
    -- CP-element group 788: 	776 
    -- CP-element group 788: successors 
    -- CP-element group 788:  members (5) 
      -- CP-element group 788: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_sample_completed_
      -- CP-element group 788: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Sample/$exit
      -- CP-element group 788: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Sample/word_access_start/$exit
      -- CP-element group 788: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Sample/word_access_start/word_0/$exit
      -- CP-element group 788: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Sample/word_access_start/word_0/ra
      -- 
    ra_10587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 788_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4820_load_0_ack_0, ack => zeropad3D_CP_2067_elements(788)); -- 
    -- CP-element group 789:  transition  input  output  bypass 
    -- CP-element group 789: predecessors 
    -- CP-element group 789: 	776 
    -- CP-element group 789: successors 
    -- CP-element group 789: 	790 
    -- CP-element group 789:  members (12) 
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_update_completed_
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/$exit
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/word_access_complete/$exit
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/word_access_complete/word_0/$exit
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/word_access_complete/word_0/ca
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/LOAD_row_high_4820_Merge/$entry
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/LOAD_row_high_4820_Merge/$exit
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/LOAD_row_high_4820_Merge/merge_req
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/LOAD_row_high_4820_Update/LOAD_row_high_4820_Merge/merge_ack
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_sample_start_
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_Sample/$entry
      -- CP-element group 789: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_Sample/rr
      -- 
    ca_10598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 789_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4820_load_0_ack_1, ack => zeropad3D_CP_2067_elements(789)); -- 
    rr_10611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(789), ack => type_cast_4824_inst_req_0); -- 
    -- CP-element group 790:  transition  input  bypass 
    -- CP-element group 790: predecessors 
    -- CP-element group 790: 	789 
    -- CP-element group 790: successors 
    -- CP-element group 790:  members (3) 
      -- CP-element group 790: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_sample_completed_
      -- CP-element group 790: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_Sample/$exit
      -- CP-element group 790: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_Sample/ra
      -- 
    ra_10612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 790_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4824_inst_ack_0, ack => zeropad3D_CP_2067_elements(790)); -- 
    -- CP-element group 791:  transition  input  bypass 
    -- CP-element group 791: predecessors 
    -- CP-element group 791: 	776 
    -- CP-element group 791: successors 
    -- CP-element group 791: 	792 
    -- CP-element group 791:  members (3) 
      -- CP-element group 791: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_update_completed_
      -- CP-element group 791: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_Update/$exit
      -- CP-element group 791: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/type_cast_4824_Update/ca
      -- 
    ca_10617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 791_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4824_inst_ack_1, ack => zeropad3D_CP_2067_elements(791)); -- 
    -- CP-element group 792:  branch  join  transition  place  output  bypass 
    -- CP-element group 792: predecessors 
    -- CP-element group 792: 	787 
    -- CP-element group 792: 	791 
    -- CP-element group 792: successors 
    -- CP-element group 792: 	793 
    -- CP-element group 792: 	794 
    -- CP-element group 792:  members (10) 
      -- CP-element group 792: 	 branch_block_stmt_655/if_stmt_4836__entry__
      -- CP-element group 792: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835__exit__
      -- CP-element group 792: 	 branch_block_stmt_655/assign_stmt_4776_to_assign_stmt_4835/$exit
      -- CP-element group 792: 	 branch_block_stmt_655/if_stmt_4836_dead_link/$entry
      -- CP-element group 792: 	 branch_block_stmt_655/if_stmt_4836_eval_test/$entry
      -- CP-element group 792: 	 branch_block_stmt_655/if_stmt_4836_eval_test/$exit
      -- CP-element group 792: 	 branch_block_stmt_655/if_stmt_4836_eval_test/branch_req
      -- CP-element group 792: 	 branch_block_stmt_655/R_cmp1696_4837_place
      -- CP-element group 792: 	 branch_block_stmt_655/if_stmt_4836_if_link/$entry
      -- CP-element group 792: 	 branch_block_stmt_655/if_stmt_4836_else_link/$entry
      -- 
    branch_req_10625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(792), ack => if_stmt_4836_branch_req_0); -- 
    zeropad3D_cp_element_group_792: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_792"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(787) & zeropad3D_CP_2067_elements(791);
      gj_zeropad3D_cp_element_group_792 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(792), clk => clk, reset => reset); --
    end block;
    -- CP-element group 793:  fork  transition  place  input  output  bypass 
    -- CP-element group 793: predecessors 
    -- CP-element group 793: 	792 
    -- CP-element group 793: successors 
    -- CP-element group 793: 	795 
    -- CP-element group 793: 	796 
    -- CP-element group 793:  members (18) 
      -- CP-element group 793: 	 branch_block_stmt_655/merge_stmt_4864__exit__
      -- CP-element group 793: 	 branch_block_stmt_655/call_stmt_4866__entry__
      -- CP-element group 793: 	 branch_block_stmt_655/if_stmt_4836_if_link/$exit
      -- CP-element group 793: 	 branch_block_stmt_655/if_stmt_4836_if_link/if_choice_transition
      -- CP-element group 793: 	 branch_block_stmt_655/ifx_xelse1670_whilex_xend1706
      -- CP-element group 793: 	 branch_block_stmt_655/call_stmt_4866/$entry
      -- CP-element group 793: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_sample_start_
      -- CP-element group 793: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_update_start_
      -- CP-element group 793: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_Sample/$entry
      -- CP-element group 793: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_Sample/crr
      -- CP-element group 793: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_Update/$entry
      -- CP-element group 793: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_Update/ccr
      -- CP-element group 793: 	 branch_block_stmt_655/ifx_xelse1670_whilex_xend1706_PhiReq/$entry
      -- CP-element group 793: 	 branch_block_stmt_655/ifx_xelse1670_whilex_xend1706_PhiReq/$exit
      -- CP-element group 793: 	 branch_block_stmt_655/merge_stmt_4864_PhiReqMerge
      -- CP-element group 793: 	 branch_block_stmt_655/merge_stmt_4864_PhiAck/$entry
      -- CP-element group 793: 	 branch_block_stmt_655/merge_stmt_4864_PhiAck/$exit
      -- CP-element group 793: 	 branch_block_stmt_655/merge_stmt_4864_PhiAck/dummy
      -- 
    if_choice_transition_10630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 793_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4836_branch_ack_1, ack => zeropad3D_CP_2067_elements(793)); -- 
    crr_10647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_10647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(793), ack => call_stmt_4866_call_req_0); -- 
    ccr_10652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_10652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(793), ack => call_stmt_4866_call_req_1); -- 
    -- CP-element group 794:  fork  transition  place  input  output  bypass 
    -- CP-element group 794: predecessors 
    -- CP-element group 794: 	792 
    -- CP-element group 794: successors 
    -- CP-element group 794: 	1228 
    -- CP-element group 794: 	1229 
    -- CP-element group 794: 	1231 
    -- CP-element group 794: 	1232 
    -- CP-element group 794: 	1233 
    -- CP-element group 794:  members (22) 
      -- CP-element group 794: 	 branch_block_stmt_655/if_stmt_4836_else_link/$exit
      -- CP-element group 794: 	 branch_block_stmt_655/if_stmt_4836_else_link/else_choice_transition
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/Sample/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/Sample/rr
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/Update/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/Update/cr
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4843/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/Sample/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/Sample/rr
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/Update/$entry
      -- CP-element group 794: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/Update/cr
      -- 
    else_choice_transition_10634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 794_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4836_branch_ack_0, ack => zeropad3D_CP_2067_elements(794)); -- 
    rr_13879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(794), ack => type_cast_4861_inst_req_0); -- 
    cr_13884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(794), ack => type_cast_4861_inst_req_1); -- 
    rr_13910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(794), ack => type_cast_4855_inst_req_0); -- 
    cr_13915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(794), ack => type_cast_4855_inst_req_1); -- 
    -- CP-element group 795:  transition  input  bypass 
    -- CP-element group 795: predecessors 
    -- CP-element group 795: 	793 
    -- CP-element group 795: successors 
    -- CP-element group 795:  members (3) 
      -- CP-element group 795: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_sample_completed_
      -- CP-element group 795: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_Sample/$exit
      -- CP-element group 795: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_Sample/cra
      -- 
    cra_10648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 795_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_4866_call_ack_0, ack => zeropad3D_CP_2067_elements(795)); -- 
    -- CP-element group 796:  transition  place  input  bypass 
    -- CP-element group 796: predecessors 
    -- CP-element group 796: 	793 
    -- CP-element group 796: successors 
    -- CP-element group 796:  members (16) 
      -- CP-element group 796: 	 branch_block_stmt_655/return__
      -- CP-element group 796: 	 branch_block_stmt_655/merge_stmt_4868__exit__
      -- CP-element group 796: 	 branch_block_stmt_655/call_stmt_4866__exit__
      -- CP-element group 796: 	 $exit
      -- CP-element group 796: 	 branch_block_stmt_655/$exit
      -- CP-element group 796: 	 branch_block_stmt_655/branch_block_stmt_655__exit__
      -- CP-element group 796: 	 branch_block_stmt_655/call_stmt_4866/$exit
      -- CP-element group 796: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_update_completed_
      -- CP-element group 796: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_Update/$exit
      -- CP-element group 796: 	 branch_block_stmt_655/call_stmt_4866/call_stmt_4866_Update/cca
      -- CP-element group 796: 	 branch_block_stmt_655/return___PhiReq/$entry
      -- CP-element group 796: 	 branch_block_stmt_655/return___PhiReq/$exit
      -- CP-element group 796: 	 branch_block_stmt_655/merge_stmt_4868_PhiReqMerge
      -- CP-element group 796: 	 branch_block_stmt_655/merge_stmt_4868_PhiAck/$entry
      -- CP-element group 796: 	 branch_block_stmt_655/merge_stmt_4868_PhiAck/$exit
      -- CP-element group 796: 	 branch_block_stmt_655/merge_stmt_4868_PhiAck/dummy
      -- 
    cca_10653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 796_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_4866_call_ack_1, ack => zeropad3D_CP_2067_elements(796)); -- 
    -- CP-element group 797:  transition  output  delay-element  bypass 
    -- CP-element group 797: predecessors 
    -- CP-element group 797: 	33 
    -- CP-element group 797: successors 
    -- CP-element group 797: 	800 
    -- CP-element group 797:  members (4) 
      -- CP-element group 797: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_747/$exit
      -- CP-element group 797: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/$exit
      -- CP-element group 797: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_751_konst_delay_trans
      -- CP-element group 797: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_req
      -- 
    phi_stmt_747_req_10664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_747_req_10664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(797), ack => phi_stmt_747_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(797) is a control-delay.
    cp_element_797_delay: control_delay_element  generic map(name => " 797_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(33), ack => zeropad3D_CP_2067_elements(797), clk => clk, reset =>reset);
    -- CP-element group 798:  transition  output  delay-element  bypass 
    -- CP-element group 798: predecessors 
    -- CP-element group 798: 	33 
    -- CP-element group 798: successors 
    -- CP-element group 798: 	800 
    -- CP-element group 798:  members (4) 
      -- CP-element group 798: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_754/$exit
      -- CP-element group 798: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/$exit
      -- CP-element group 798: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_758_konst_delay_trans
      -- CP-element group 798: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_req
      -- 
    phi_stmt_754_req_10672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_754_req_10672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(798), ack => phi_stmt_754_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(798) is a control-delay.
    cp_element_798_delay: control_delay_element  generic map(name => " 798_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(33), ack => zeropad3D_CP_2067_elements(798), clk => clk, reset =>reset);
    -- CP-element group 799:  transition  output  delay-element  bypass 
    -- CP-element group 799: predecessors 
    -- CP-element group 799: 	33 
    -- CP-element group 799: successors 
    -- CP-element group 799: 	800 
    -- CP-element group 799:  members (4) 
      -- CP-element group 799: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_761/$exit
      -- CP-element group 799: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/$exit
      -- CP-element group 799: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_765_konst_delay_trans
      -- CP-element group 799: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_req
      -- 
    phi_stmt_761_req_10680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_761_req_10680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(799), ack => phi_stmt_761_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(799) is a control-delay.
    cp_element_799_delay: control_delay_element  generic map(name => " 799_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(33), ack => zeropad3D_CP_2067_elements(799), clk => clk, reset =>reset);
    -- CP-element group 800:  join  transition  bypass 
    -- CP-element group 800: predecessors 
    -- CP-element group 800: 	797 
    -- CP-element group 800: 	798 
    -- CP-element group 800: 	799 
    -- CP-element group 800: successors 
    -- CP-element group 800: 	811 
    -- CP-element group 800:  members (1) 
      -- CP-element group 800: 	 branch_block_stmt_655/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_800: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_800"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(797) & zeropad3D_CP_2067_elements(798) & zeropad3D_CP_2067_elements(799);
      gj_zeropad3D_cp_element_group_800 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(800), clk => clk, reset => reset); --
    end block;
    -- CP-element group 801:  transition  input  bypass 
    -- CP-element group 801: predecessors 
    -- CP-element group 801: 	1 
    -- CP-element group 801: successors 
    -- CP-element group 801: 	803 
    -- CP-element group 801:  members (2) 
      -- CP-element group 801: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/Sample/$exit
      -- CP-element group 801: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/Sample/ra
      -- 
    ra_10700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 801_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_753_inst_ack_0, ack => zeropad3D_CP_2067_elements(801)); -- 
    -- CP-element group 802:  transition  input  bypass 
    -- CP-element group 802: predecessors 
    -- CP-element group 802: 	1 
    -- CP-element group 802: successors 
    -- CP-element group 802: 	803 
    -- CP-element group 802:  members (2) 
      -- CP-element group 802: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/Update/$exit
      -- CP-element group 802: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/Update/ca
      -- 
    ca_10705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 802_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_753_inst_ack_1, ack => zeropad3D_CP_2067_elements(802)); -- 
    -- CP-element group 803:  join  transition  output  bypass 
    -- CP-element group 803: predecessors 
    -- CP-element group 803: 	801 
    -- CP-element group 803: 	802 
    -- CP-element group 803: successors 
    -- CP-element group 803: 	810 
    -- CP-element group 803:  members (5) 
      -- CP-element group 803: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/$exit
      -- CP-element group 803: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/$exit
      -- CP-element group 803: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/$exit
      -- CP-element group 803: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_sources/type_cast_753/SplitProtocol/$exit
      -- CP-element group 803: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_747/phi_stmt_747_req
      -- 
    phi_stmt_747_req_10706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_747_req_10706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(803), ack => phi_stmt_747_req_1); -- 
    zeropad3D_cp_element_group_803: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_803"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(801) & zeropad3D_CP_2067_elements(802);
      gj_zeropad3D_cp_element_group_803 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(803), clk => clk, reset => reset); --
    end block;
    -- CP-element group 804:  transition  input  bypass 
    -- CP-element group 804: predecessors 
    -- CP-element group 804: 	1 
    -- CP-element group 804: successors 
    -- CP-element group 804: 	806 
    -- CP-element group 804:  members (2) 
      -- CP-element group 804: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/Sample/$exit
      -- CP-element group 804: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/Sample/ra
      -- 
    ra_10723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 804_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_760_inst_ack_0, ack => zeropad3D_CP_2067_elements(804)); -- 
    -- CP-element group 805:  transition  input  bypass 
    -- CP-element group 805: predecessors 
    -- CP-element group 805: 	1 
    -- CP-element group 805: successors 
    -- CP-element group 805: 	806 
    -- CP-element group 805:  members (2) 
      -- CP-element group 805: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/Update/$exit
      -- CP-element group 805: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/Update/ca
      -- 
    ca_10728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 805_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_760_inst_ack_1, ack => zeropad3D_CP_2067_elements(805)); -- 
    -- CP-element group 806:  join  transition  output  bypass 
    -- CP-element group 806: predecessors 
    -- CP-element group 806: 	804 
    -- CP-element group 806: 	805 
    -- CP-element group 806: successors 
    -- CP-element group 806: 	810 
    -- CP-element group 806:  members (5) 
      -- CP-element group 806: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/$exit
      -- CP-element group 806: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/$exit
      -- CP-element group 806: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/$exit
      -- CP-element group 806: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_sources/type_cast_760/SplitProtocol/$exit
      -- CP-element group 806: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_754/phi_stmt_754_req
      -- 
    phi_stmt_754_req_10729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_754_req_10729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(806), ack => phi_stmt_754_req_1); -- 
    zeropad3D_cp_element_group_806: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_806"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(804) & zeropad3D_CP_2067_elements(805);
      gj_zeropad3D_cp_element_group_806 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(806), clk => clk, reset => reset); --
    end block;
    -- CP-element group 807:  transition  input  bypass 
    -- CP-element group 807: predecessors 
    -- CP-element group 807: 	1 
    -- CP-element group 807: successors 
    -- CP-element group 807: 	809 
    -- CP-element group 807:  members (2) 
      -- CP-element group 807: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/Sample/$exit
      -- CP-element group 807: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/Sample/ra
      -- 
    ra_10746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 807_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_767_inst_ack_0, ack => zeropad3D_CP_2067_elements(807)); -- 
    -- CP-element group 808:  transition  input  bypass 
    -- CP-element group 808: predecessors 
    -- CP-element group 808: 	1 
    -- CP-element group 808: successors 
    -- CP-element group 808: 	809 
    -- CP-element group 808:  members (2) 
      -- CP-element group 808: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/Update/$exit
      -- CP-element group 808: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/Update/ca
      -- 
    ca_10751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 808_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_767_inst_ack_1, ack => zeropad3D_CP_2067_elements(808)); -- 
    -- CP-element group 809:  join  transition  output  bypass 
    -- CP-element group 809: predecessors 
    -- CP-element group 809: 	807 
    -- CP-element group 809: 	808 
    -- CP-element group 809: successors 
    -- CP-element group 809: 	810 
    -- CP-element group 809:  members (5) 
      -- CP-element group 809: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/$exit
      -- CP-element group 809: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/$exit
      -- CP-element group 809: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/$exit
      -- CP-element group 809: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_sources/type_cast_767/SplitProtocol/$exit
      -- CP-element group 809: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/phi_stmt_761/phi_stmt_761_req
      -- 
    phi_stmt_761_req_10752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_761_req_10752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(809), ack => phi_stmt_761_req_1); -- 
    zeropad3D_cp_element_group_809: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_809"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(807) & zeropad3D_CP_2067_elements(808);
      gj_zeropad3D_cp_element_group_809 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(809), clk => clk, reset => reset); --
    end block;
    -- CP-element group 810:  join  transition  bypass 
    -- CP-element group 810: predecessors 
    -- CP-element group 810: 	803 
    -- CP-element group 810: 	806 
    -- CP-element group 810: 	809 
    -- CP-element group 810: successors 
    -- CP-element group 810: 	811 
    -- CP-element group 810:  members (1) 
      -- CP-element group 810: 	 branch_block_stmt_655/ifx_xend174_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_810: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_810"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(803) & zeropad3D_CP_2067_elements(806) & zeropad3D_CP_2067_elements(809);
      gj_zeropad3D_cp_element_group_810 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(810), clk => clk, reset => reset); --
    end block;
    -- CP-element group 811:  merge  fork  transition  place  bypass 
    -- CP-element group 811: predecessors 
    -- CP-element group 811: 	800 
    -- CP-element group 811: 	810 
    -- CP-element group 811: successors 
    -- CP-element group 811: 	812 
    -- CP-element group 811: 	813 
    -- CP-element group 811: 	814 
    -- CP-element group 811:  members (2) 
      -- CP-element group 811: 	 branch_block_stmt_655/merge_stmt_746_PhiReqMerge
      -- CP-element group 811: 	 branch_block_stmt_655/merge_stmt_746_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(811) <= OrReduce(zeropad3D_CP_2067_elements(800) & zeropad3D_CP_2067_elements(810));
    -- CP-element group 812:  transition  input  bypass 
    -- CP-element group 812: predecessors 
    -- CP-element group 812: 	811 
    -- CP-element group 812: successors 
    -- CP-element group 812: 	815 
    -- CP-element group 812:  members (1) 
      -- CP-element group 812: 	 branch_block_stmt_655/merge_stmt_746_PhiAck/phi_stmt_747_ack
      -- 
    phi_stmt_747_ack_10757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 812_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_747_ack_0, ack => zeropad3D_CP_2067_elements(812)); -- 
    -- CP-element group 813:  transition  input  bypass 
    -- CP-element group 813: predecessors 
    -- CP-element group 813: 	811 
    -- CP-element group 813: successors 
    -- CP-element group 813: 	815 
    -- CP-element group 813:  members (1) 
      -- CP-element group 813: 	 branch_block_stmt_655/merge_stmt_746_PhiAck/phi_stmt_754_ack
      -- 
    phi_stmt_754_ack_10758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 813_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_754_ack_0, ack => zeropad3D_CP_2067_elements(813)); -- 
    -- CP-element group 814:  transition  input  bypass 
    -- CP-element group 814: predecessors 
    -- CP-element group 814: 	811 
    -- CP-element group 814: successors 
    -- CP-element group 814: 	815 
    -- CP-element group 814:  members (1) 
      -- CP-element group 814: 	 branch_block_stmt_655/merge_stmt_746_PhiAck/phi_stmt_761_ack
      -- 
    phi_stmt_761_ack_10759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 814_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_761_ack_0, ack => zeropad3D_CP_2067_elements(814)); -- 
    -- CP-element group 815:  join  fork  transition  place  output  bypass 
    -- CP-element group 815: predecessors 
    -- CP-element group 815: 	812 
    -- CP-element group 815: 	813 
    -- CP-element group 815: 	814 
    -- CP-element group 815: successors 
    -- CP-element group 815: 	34 
    -- CP-element group 815: 	35 
    -- CP-element group 815:  members (10) 
      -- CP-element group 815: 	 branch_block_stmt_655/merge_stmt_746__exit__
      -- CP-element group 815: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780__entry__
      -- CP-element group 815: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/$entry
      -- CP-element group 815: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_sample_start_
      -- CP-element group 815: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_update_start_
      -- CP-element group 815: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_Sample/$entry
      -- CP-element group 815: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_Sample/rr
      -- CP-element group 815: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_Update/$entry
      -- CP-element group 815: 	 branch_block_stmt_655/assign_stmt_773_to_assign_stmt_780/type_cast_772_Update/cr
      -- CP-element group 815: 	 branch_block_stmt_655/merge_stmt_746_PhiAck/$exit
      -- 
    rr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(815), ack => type_cast_772_inst_req_0); -- 
    cr_2797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(815), ack => type_cast_772_inst_req_1); -- 
    zeropad3D_cp_element_group_815: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_815"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(812) & zeropad3D_CP_2067_elements(813) & zeropad3D_CP_2067_elements(814);
      gj_zeropad3D_cp_element_group_815 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(815), clk => clk, reset => reset); --
    end block;
    -- CP-element group 816:  merge  fork  transition  place  output  bypass 
    -- CP-element group 816: predecessors 
    -- CP-element group 816: 	36 
    -- CP-element group 816: 	43 
    -- CP-element group 816: 	46 
    -- CP-element group 816: 	53 
    -- CP-element group 816: successors 
    -- CP-element group 816: 	56 
    -- CP-element group 816: 	57 
    -- CP-element group 816: 	60 
    -- CP-element group 816: 	62 
    -- CP-element group 816: 	64 
    -- CP-element group 816: 	66 
    -- CP-element group 816: 	54 
    -- CP-element group 816: 	55 
    -- CP-element group 816:  members (33) 
      -- CP-element group 816: 	 branch_block_stmt_655/merge_stmt_870__exit__
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927__entry__
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_sample_start_
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_update_start_
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_Sample/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_Sample/rr
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_Update/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_874_Update/cr
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_sample_start_
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_update_start_
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_Sample/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_Sample/rr
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_Update/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_879_Update/cr
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_update_start_
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_Update/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/type_cast_914_Update/cr
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_update_start_
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_update_start
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_Update/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/array_obj_ref_920_final_index_sum_regn_Update/req
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_complete/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/addr_of_921_complete/req
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_update_start_
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Update/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Update/word_access_complete/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Update/word_access_complete/word_0/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/assign_stmt_875_to_assign_stmt_927/ptr_deref_924_Update/word_access_complete/word_0/cr
      -- CP-element group 816: 	 branch_block_stmt_655/merge_stmt_870_PhiReqMerge
      -- CP-element group 816: 	 branch_block_stmt_655/merge_stmt_870_PhiAck/$entry
      -- CP-element group 816: 	 branch_block_stmt_655/merge_stmt_870_PhiAck/$exit
      -- CP-element group 816: 	 branch_block_stmt_655/merge_stmt_870_PhiAck/dummy
      -- 
    rr_3002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(816), ack => type_cast_874_inst_req_0); -- 
    cr_3007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(816), ack => type_cast_874_inst_req_1); -- 
    rr_3016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(816), ack => type_cast_879_inst_req_0); -- 
    cr_3021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(816), ack => type_cast_879_inst_req_1); -- 
    cr_3035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(816), ack => type_cast_914_inst_req_1); -- 
    req_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(816), ack => array_obj_ref_920_index_offset_req_1); -- 
    req_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(816), ack => addr_of_921_final_reg_req_1); -- 
    cr_3131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(816), ack => ptr_deref_924_store_0_req_1); -- 
    zeropad3D_CP_2067_elements(816) <= OrReduce(zeropad3D_CP_2067_elements(36) & zeropad3D_CP_2067_elements(43) & zeropad3D_CP_2067_elements(46) & zeropad3D_CP_2067_elements(53));
    -- CP-element group 817:  merge  fork  transition  place  output  bypass 
    -- CP-element group 817: predecessors 
    -- CP-element group 817: 	67 
    -- CP-element group 817: 	87 
    -- CP-element group 817: successors 
    -- CP-element group 817: 	88 
    -- CP-element group 817: 	89 
    -- CP-element group 817:  members (13) 
      -- CP-element group 817: 	 branch_block_stmt_655/merge_stmt_1036__exit__
      -- CP-element group 817: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054__entry__
      -- CP-element group 817: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/$entry
      -- CP-element group 817: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_sample_start_
      -- CP-element group 817: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_update_start_
      -- CP-element group 817: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_Sample/$entry
      -- CP-element group 817: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_Sample/rr
      -- CP-element group 817: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_Update/$entry
      -- CP-element group 817: 	 branch_block_stmt_655/assign_stmt_1041_to_assign_stmt_1054/type_cast_1040_Update/cr
      -- CP-element group 817: 	 branch_block_stmt_655/merge_stmt_1036_PhiReqMerge
      -- CP-element group 817: 	 branch_block_stmt_655/merge_stmt_1036_PhiAck/$entry
      -- CP-element group 817: 	 branch_block_stmt_655/merge_stmt_1036_PhiAck/$exit
      -- CP-element group 817: 	 branch_block_stmt_655/merge_stmt_1036_PhiAck/dummy
      -- 
    rr_3380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(817), ack => type_cast_1040_inst_req_0); -- 
    cr_3385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(817), ack => type_cast_1040_inst_req_1); -- 
    zeropad3D_CP_2067_elements(817) <= OrReduce(zeropad3D_CP_2067_elements(67) & zeropad3D_CP_2067_elements(87));
    -- CP-element group 818:  transition  input  bypass 
    -- CP-element group 818: predecessors 
    -- CP-element group 818: 	109 
    -- CP-element group 818: successors 
    -- CP-element group 818: 	820 
    -- CP-element group 818:  members (2) 
      -- CP-element group 818: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/Sample/$exit
      -- CP-element group 818: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/Sample/ra
      -- 
    ra_10879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 818_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_0, ack => zeropad3D_CP_2067_elements(818)); -- 
    -- CP-element group 819:  transition  input  bypass 
    -- CP-element group 819: predecessors 
    -- CP-element group 819: 	109 
    -- CP-element group 819: successors 
    -- CP-element group 819: 	820 
    -- CP-element group 819:  members (2) 
      -- CP-element group 819: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/Update/$exit
      -- CP-element group 819: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/Update/ca
      -- 
    ca_10884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 819_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_1, ack => zeropad3D_CP_2067_elements(819)); -- 
    -- CP-element group 820:  join  transition  output  bypass 
    -- CP-element group 820: predecessors 
    -- CP-element group 820: 	818 
    -- CP-element group 820: 	819 
    -- CP-element group 820: successors 
    -- CP-element group 820: 	825 
    -- CP-element group 820:  members (5) 
      -- CP-element group 820: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/$exit
      -- CP-element group 820: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/$exit
      -- CP-element group 820: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/$exit
      -- CP-element group 820: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1160/SplitProtocol/$exit
      -- CP-element group 820: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_req
      -- 
    phi_stmt_1155_req_10885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1155_req_10885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(820), ack => phi_stmt_1155_req_1); -- 
    zeropad3D_cp_element_group_820: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_820"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(818) & zeropad3D_CP_2067_elements(819);
      gj_zeropad3D_cp_element_group_820 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(820), clk => clk, reset => reset); --
    end block;
    -- CP-element group 821:  transition  input  bypass 
    -- CP-element group 821: predecessors 
    -- CP-element group 821: 	109 
    -- CP-element group 821: successors 
    -- CP-element group 821: 	823 
    -- CP-element group 821:  members (2) 
      -- CP-element group 821: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/Sample/$exit
      -- CP-element group 821: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/Sample/ra
      -- 
    ra_10902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 821_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1166_inst_ack_0, ack => zeropad3D_CP_2067_elements(821)); -- 
    -- CP-element group 822:  transition  input  bypass 
    -- CP-element group 822: predecessors 
    -- CP-element group 822: 	109 
    -- CP-element group 822: successors 
    -- CP-element group 822: 	823 
    -- CP-element group 822:  members (2) 
      -- CP-element group 822: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/Update/$exit
      -- CP-element group 822: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/Update/ca
      -- 
    ca_10907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 822_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1166_inst_ack_1, ack => zeropad3D_CP_2067_elements(822)); -- 
    -- CP-element group 823:  join  transition  output  bypass 
    -- CP-element group 823: predecessors 
    -- CP-element group 823: 	821 
    -- CP-element group 823: 	822 
    -- CP-element group 823: successors 
    -- CP-element group 823: 	825 
    -- CP-element group 823:  members (5) 
      -- CP-element group 823: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/$exit
      -- CP-element group 823: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/$exit
      -- CP-element group 823: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/$exit
      -- CP-element group 823: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1166/SplitProtocol/$exit
      -- CP-element group 823: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_req
      -- 
    phi_stmt_1161_req_10908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1161_req_10908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(823), ack => phi_stmt_1161_req_1); -- 
    zeropad3D_cp_element_group_823: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_823"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(821) & zeropad3D_CP_2067_elements(822);
      gj_zeropad3D_cp_element_group_823 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(823), clk => clk, reset => reset); --
    end block;
    -- CP-element group 824:  transition  output  delay-element  bypass 
    -- CP-element group 824: predecessors 
    -- CP-element group 824: 	109 
    -- CP-element group 824: successors 
    -- CP-element group 824: 	825 
    -- CP-element group 824:  members (4) 
      -- CP-element group 824: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1167/$exit
      -- CP-element group 824: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/$exit
      -- CP-element group 824: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1173_konst_delay_trans
      -- CP-element group 824: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_req
      -- 
    phi_stmt_1167_req_10916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1167_req_10916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(824), ack => phi_stmt_1167_req_1); -- 
    -- Element group zeropad3D_CP_2067_elements(824) is a control-delay.
    cp_element_824_delay: control_delay_element  generic map(name => " 824_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(109), ack => zeropad3D_CP_2067_elements(824), clk => clk, reset =>reset);
    -- CP-element group 825:  join  transition  bypass 
    -- CP-element group 825: predecessors 
    -- CP-element group 825: 	820 
    -- CP-element group 825: 	823 
    -- CP-element group 825: 	824 
    -- CP-element group 825: successors 
    -- CP-element group 825: 	836 
    -- CP-element group 825:  members (1) 
      -- CP-element group 825: 	 branch_block_stmt_655/ifx_xelse140_ifx_xend174_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_825: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_825"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(820) & zeropad3D_CP_2067_elements(823) & zeropad3D_CP_2067_elements(824);
      gj_zeropad3D_cp_element_group_825 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(825), clk => clk, reset => reset); --
    end block;
    -- CP-element group 826:  transition  input  bypass 
    -- CP-element group 826: predecessors 
    -- CP-element group 826: 	90 
    -- CP-element group 826: successors 
    -- CP-element group 826: 	828 
    -- CP-element group 826:  members (2) 
      -- CP-element group 826: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/Sample/$exit
      -- CP-element group 826: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/Sample/ra
      -- 
    ra_10936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 826_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1158_inst_ack_0, ack => zeropad3D_CP_2067_elements(826)); -- 
    -- CP-element group 827:  transition  input  bypass 
    -- CP-element group 827: predecessors 
    -- CP-element group 827: 	90 
    -- CP-element group 827: successors 
    -- CP-element group 827: 	828 
    -- CP-element group 827:  members (2) 
      -- CP-element group 827: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/Update/$exit
      -- CP-element group 827: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/Update/ca
      -- 
    ca_10941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 827_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1158_inst_ack_1, ack => zeropad3D_CP_2067_elements(827)); -- 
    -- CP-element group 828:  join  transition  output  bypass 
    -- CP-element group 828: predecessors 
    -- CP-element group 828: 	826 
    -- CP-element group 828: 	827 
    -- CP-element group 828: successors 
    -- CP-element group 828: 	835 
    -- CP-element group 828:  members (5) 
      -- CP-element group 828: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/$exit
      -- CP-element group 828: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/$exit
      -- CP-element group 828: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/$exit
      -- CP-element group 828: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_sources/type_cast_1158/SplitProtocol/$exit
      -- CP-element group 828: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1155/phi_stmt_1155_req
      -- 
    phi_stmt_1155_req_10942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1155_req_10942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(828), ack => phi_stmt_1155_req_0); -- 
    zeropad3D_cp_element_group_828: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_828"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(826) & zeropad3D_CP_2067_elements(827);
      gj_zeropad3D_cp_element_group_828 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(828), clk => clk, reset => reset); --
    end block;
    -- CP-element group 829:  transition  input  bypass 
    -- CP-element group 829: predecessors 
    -- CP-element group 829: 	90 
    -- CP-element group 829: successors 
    -- CP-element group 829: 	831 
    -- CP-element group 829:  members (2) 
      -- CP-element group 829: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Sample/$exit
      -- CP-element group 829: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Sample/ra
      -- 
    ra_10959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 829_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1164_inst_ack_0, ack => zeropad3D_CP_2067_elements(829)); -- 
    -- CP-element group 830:  transition  input  bypass 
    -- CP-element group 830: predecessors 
    -- CP-element group 830: 	90 
    -- CP-element group 830: successors 
    -- CP-element group 830: 	831 
    -- CP-element group 830:  members (2) 
      -- CP-element group 830: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Update/$exit
      -- CP-element group 830: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Update/ca
      -- 
    ca_10964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 830_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1164_inst_ack_1, ack => zeropad3D_CP_2067_elements(830)); -- 
    -- CP-element group 831:  join  transition  output  bypass 
    -- CP-element group 831: predecessors 
    -- CP-element group 831: 	829 
    -- CP-element group 831: 	830 
    -- CP-element group 831: successors 
    -- CP-element group 831: 	835 
    -- CP-element group 831:  members (5) 
      -- CP-element group 831: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/$exit
      -- CP-element group 831: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/$exit
      -- CP-element group 831: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/$exit
      -- CP-element group 831: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/$exit
      -- CP-element group 831: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1161/phi_stmt_1161_req
      -- 
    phi_stmt_1161_req_10965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1161_req_10965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(831), ack => phi_stmt_1161_req_0); -- 
    zeropad3D_cp_element_group_831: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_831"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(829) & zeropad3D_CP_2067_elements(830);
      gj_zeropad3D_cp_element_group_831 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(831), clk => clk, reset => reset); --
    end block;
    -- CP-element group 832:  transition  input  bypass 
    -- CP-element group 832: predecessors 
    -- CP-element group 832: 	90 
    -- CP-element group 832: successors 
    -- CP-element group 832: 	834 
    -- CP-element group 832:  members (2) 
      -- CP-element group 832: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/Sample/$exit
      -- CP-element group 832: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/Sample/ra
      -- 
    ra_10982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 832_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1170_inst_ack_0, ack => zeropad3D_CP_2067_elements(832)); -- 
    -- CP-element group 833:  transition  input  bypass 
    -- CP-element group 833: predecessors 
    -- CP-element group 833: 	90 
    -- CP-element group 833: successors 
    -- CP-element group 833: 	834 
    -- CP-element group 833:  members (2) 
      -- CP-element group 833: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/Update/$exit
      -- CP-element group 833: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/Update/ca
      -- 
    ca_10987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 833_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1170_inst_ack_1, ack => zeropad3D_CP_2067_elements(833)); -- 
    -- CP-element group 834:  join  transition  output  bypass 
    -- CP-element group 834: predecessors 
    -- CP-element group 834: 	832 
    -- CP-element group 834: 	833 
    -- CP-element group 834: successors 
    -- CP-element group 834: 	835 
    -- CP-element group 834:  members (5) 
      -- CP-element group 834: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/$exit
      -- CP-element group 834: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/$exit
      -- CP-element group 834: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/$exit
      -- CP-element group 834: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_sources/type_cast_1170/SplitProtocol/$exit
      -- CP-element group 834: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/phi_stmt_1167/phi_stmt_1167_req
      -- 
    phi_stmt_1167_req_10988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1167_req_10988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(834), ack => phi_stmt_1167_req_0); -- 
    zeropad3D_cp_element_group_834: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_834"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(832) & zeropad3D_CP_2067_elements(833);
      gj_zeropad3D_cp_element_group_834 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(834), clk => clk, reset => reset); --
    end block;
    -- CP-element group 835:  join  transition  bypass 
    -- CP-element group 835: predecessors 
    -- CP-element group 835: 	828 
    -- CP-element group 835: 	831 
    -- CP-element group 835: 	834 
    -- CP-element group 835: successors 
    -- CP-element group 835: 	836 
    -- CP-element group 835:  members (1) 
      -- CP-element group 835: 	 branch_block_stmt_655/ifx_xthen135_ifx_xend174_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_835: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_835"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(828) & zeropad3D_CP_2067_elements(831) & zeropad3D_CP_2067_elements(834);
      gj_zeropad3D_cp_element_group_835 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(835), clk => clk, reset => reset); --
    end block;
    -- CP-element group 836:  merge  fork  transition  place  bypass 
    -- CP-element group 836: predecessors 
    -- CP-element group 836: 	825 
    -- CP-element group 836: 	835 
    -- CP-element group 836: successors 
    -- CP-element group 836: 	837 
    -- CP-element group 836: 	838 
    -- CP-element group 836: 	839 
    -- CP-element group 836:  members (2) 
      -- CP-element group 836: 	 branch_block_stmt_655/merge_stmt_1154_PhiReqMerge
      -- CP-element group 836: 	 branch_block_stmt_655/merge_stmt_1154_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(836) <= OrReduce(zeropad3D_CP_2067_elements(825) & zeropad3D_CP_2067_elements(835));
    -- CP-element group 837:  transition  input  bypass 
    -- CP-element group 837: predecessors 
    -- CP-element group 837: 	836 
    -- CP-element group 837: successors 
    -- CP-element group 837: 	840 
    -- CP-element group 837:  members (1) 
      -- CP-element group 837: 	 branch_block_stmt_655/merge_stmt_1154_PhiAck/phi_stmt_1155_ack
      -- 
    phi_stmt_1155_ack_10993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 837_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1155_ack_0, ack => zeropad3D_CP_2067_elements(837)); -- 
    -- CP-element group 838:  transition  input  bypass 
    -- CP-element group 838: predecessors 
    -- CP-element group 838: 	836 
    -- CP-element group 838: successors 
    -- CP-element group 838: 	840 
    -- CP-element group 838:  members (1) 
      -- CP-element group 838: 	 branch_block_stmt_655/merge_stmt_1154_PhiAck/phi_stmt_1161_ack
      -- 
    phi_stmt_1161_ack_10994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 838_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1161_ack_0, ack => zeropad3D_CP_2067_elements(838)); -- 
    -- CP-element group 839:  transition  input  bypass 
    -- CP-element group 839: predecessors 
    -- CP-element group 839: 	836 
    -- CP-element group 839: successors 
    -- CP-element group 839: 	840 
    -- CP-element group 839:  members (1) 
      -- CP-element group 839: 	 branch_block_stmt_655/merge_stmt_1154_PhiAck/phi_stmt_1167_ack
      -- 
    phi_stmt_1167_ack_10995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 839_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1167_ack_0, ack => zeropad3D_CP_2067_elements(839)); -- 
    -- CP-element group 840:  join  transition  bypass 
    -- CP-element group 840: predecessors 
    -- CP-element group 840: 	837 
    -- CP-element group 840: 	838 
    -- CP-element group 840: 	839 
    -- CP-element group 840: successors 
    -- CP-element group 840: 	1 
    -- CP-element group 840:  members (1) 
      -- CP-element group 840: 	 branch_block_stmt_655/merge_stmt_1154_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_840: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_840"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(837) & zeropad3D_CP_2067_elements(838) & zeropad3D_CP_2067_elements(839);
      gj_zeropad3D_cp_element_group_840 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(840), clk => clk, reset => reset); --
    end block;
    -- CP-element group 841:  transition  input  bypass 
    -- CP-element group 841: predecessors 
    -- CP-element group 841: 	108 
    -- CP-element group 841: successors 
    -- CP-element group 841: 	843 
    -- CP-element group 841:  members (2) 
      -- CP-element group 841: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/Sample/$exit
      -- CP-element group 841: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/Sample/ra
      -- 
    ra_11015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 841_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1180_inst_ack_0, ack => zeropad3D_CP_2067_elements(841)); -- 
    -- CP-element group 842:  transition  input  bypass 
    -- CP-element group 842: predecessors 
    -- CP-element group 842: 	108 
    -- CP-element group 842: successors 
    -- CP-element group 842: 	843 
    -- CP-element group 842:  members (2) 
      -- CP-element group 842: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/Update/$exit
      -- CP-element group 842: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/Update/ca
      -- 
    ca_11020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 842_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1180_inst_ack_1, ack => zeropad3D_CP_2067_elements(842)); -- 
    -- CP-element group 843:  join  transition  output  bypass 
    -- CP-element group 843: predecessors 
    -- CP-element group 843: 	841 
    -- CP-element group 843: 	842 
    -- CP-element group 843: successors 
    -- CP-element group 843: 	847 
    -- CP-element group 843:  members (5) 
      -- CP-element group 843: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/$exit
      -- CP-element group 843: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/$exit
      -- CP-element group 843: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/$exit
      -- CP-element group 843: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_sources/type_cast_1180/SplitProtocol/$exit
      -- CP-element group 843: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1177/phi_stmt_1177_req
      -- 
    phi_stmt_1177_req_11021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1177_req_11021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(843), ack => phi_stmt_1177_req_0); -- 
    zeropad3D_cp_element_group_843: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_843"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(841) & zeropad3D_CP_2067_elements(842);
      gj_zeropad3D_cp_element_group_843 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(843), clk => clk, reset => reset); --
    end block;
    -- CP-element group 844:  transition  input  bypass 
    -- CP-element group 844: predecessors 
    -- CP-element group 844: 	108 
    -- CP-element group 844: successors 
    -- CP-element group 844: 	846 
    -- CP-element group 844:  members (2) 
      -- CP-element group 844: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/Sample/$exit
      -- CP-element group 844: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/Sample/ra
      -- 
    ra_11038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 844_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1184_inst_ack_0, ack => zeropad3D_CP_2067_elements(844)); -- 
    -- CP-element group 845:  transition  input  bypass 
    -- CP-element group 845: predecessors 
    -- CP-element group 845: 	108 
    -- CP-element group 845: successors 
    -- CP-element group 845: 	846 
    -- CP-element group 845:  members (2) 
      -- CP-element group 845: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/Update/$exit
      -- CP-element group 845: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/Update/ca
      -- 
    ca_11043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 845_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1184_inst_ack_1, ack => zeropad3D_CP_2067_elements(845)); -- 
    -- CP-element group 846:  join  transition  output  bypass 
    -- CP-element group 846: predecessors 
    -- CP-element group 846: 	844 
    -- CP-element group 846: 	845 
    -- CP-element group 846: successors 
    -- CP-element group 846: 	847 
    -- CP-element group 846:  members (5) 
      -- CP-element group 846: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/$exit
      -- CP-element group 846: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/$exit
      -- CP-element group 846: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/$exit
      -- CP-element group 846: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_sources/type_cast_1184/SplitProtocol/$exit
      -- CP-element group 846: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/phi_stmt_1181/phi_stmt_1181_req
      -- 
    phi_stmt_1181_req_11044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1181_req_11044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(846), ack => phi_stmt_1181_req_0); -- 
    zeropad3D_cp_element_group_846: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_846"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(844) & zeropad3D_CP_2067_elements(845);
      gj_zeropad3D_cp_element_group_846 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(846), clk => clk, reset => reset); --
    end block;
    -- CP-element group 847:  join  fork  transition  place  bypass 
    -- CP-element group 847: predecessors 
    -- CP-element group 847: 	843 
    -- CP-element group 847: 	846 
    -- CP-element group 847: successors 
    -- CP-element group 847: 	848 
    -- CP-element group 847: 	849 
    -- CP-element group 847:  members (3) 
      -- CP-element group 847: 	 branch_block_stmt_655/ifx_xelse140_whilex_xend_PhiReq/$exit
      -- CP-element group 847: 	 branch_block_stmt_655/merge_stmt_1176_PhiReqMerge
      -- CP-element group 847: 	 branch_block_stmt_655/merge_stmt_1176_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_847: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_847"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(843) & zeropad3D_CP_2067_elements(846);
      gj_zeropad3D_cp_element_group_847 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(847), clk => clk, reset => reset); --
    end block;
    -- CP-element group 848:  transition  input  bypass 
    -- CP-element group 848: predecessors 
    -- CP-element group 848: 	847 
    -- CP-element group 848: successors 
    -- CP-element group 848: 	850 
    -- CP-element group 848:  members (1) 
      -- CP-element group 848: 	 branch_block_stmt_655/merge_stmt_1176_PhiAck/phi_stmt_1177_ack
      -- 
    phi_stmt_1177_ack_11049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 848_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1177_ack_0, ack => zeropad3D_CP_2067_elements(848)); -- 
    -- CP-element group 849:  transition  input  bypass 
    -- CP-element group 849: predecessors 
    -- CP-element group 849: 	847 
    -- CP-element group 849: successors 
    -- CP-element group 849: 	850 
    -- CP-element group 849:  members (1) 
      -- CP-element group 849: 	 branch_block_stmt_655/merge_stmt_1176_PhiAck/phi_stmt_1181_ack
      -- 
    phi_stmt_1181_ack_11050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 849_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1181_ack_0, ack => zeropad3D_CP_2067_elements(849)); -- 
    -- CP-element group 850:  join  fork  transition  place  output  bypass 
    -- CP-element group 850: predecessors 
    -- CP-element group 850: 	848 
    -- CP-element group 850: 	849 
    -- CP-element group 850: successors 
    -- CP-element group 850: 	110 
    -- CP-element group 850: 	111 
    -- CP-element group 850: 	112 
    -- CP-element group 850: 	113 
    -- CP-element group 850: 	114 
    -- CP-element group 850: 	115 
    -- CP-element group 850: 	116 
    -- CP-element group 850: 	117 
    -- CP-element group 850: 	118 
    -- CP-element group 850: 	119 
    -- CP-element group 850: 	121 
    -- CP-element group 850: 	123 
    -- CP-element group 850: 	125 
    -- CP-element group 850: 	127 
    -- CP-element group 850: 	129 
    -- CP-element group 850:  members (73) 
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Sample/word_access_start/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Sample/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_root_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_word_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_root_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_Sample/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Sample/word_access_start/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_word_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_sample_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Sample/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/merge_stmt_1176__exit__
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273__entry__
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/word_access_complete/word_0/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_Update/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/word_access_complete/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/word_access_complete/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_sample_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1231_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/word_access_complete/word_0/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/word_access_complete/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Sample/word_access_start/word_0/rr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_sample_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Sample/word_access_start/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_Update/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Sample/word_access_start/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_Sample/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_root_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_word_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/word_access_complete/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_depth_high_1200_sample_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_depth_high_1203_Sample/word_access_start/word_0/rr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1227_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/word_access_complete/word_0/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/word_access_complete/word_0/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/word_access_complete/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1214_Update/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/word_access_complete/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/word_access_complete/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Sample/word_access_start/word_0/rr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Sample/word_access_start/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Sample/word_access_start/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/word_access_complete/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Sample/word_access_start/word_0/rr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1218_Update/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1210_Update/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_Sample/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_root_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_word_address_calculated
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_update_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_pad_1197_sample_start_
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Sample/word_access_start/word_0/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_Update/cr
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_Update/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/LOAD_out_col_high_1206_Sample/word_access_start/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/$entry
      -- CP-element group 850: 	 branch_block_stmt_655/assign_stmt_1189_to_assign_stmt_1273/type_cast_1188_Sample/rr
      -- CP-element group 850: 	 branch_block_stmt_655/merge_stmt_1176_PhiAck/$exit
      -- 
    cr_3643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => LOAD_depth_high_1200_load_0_req_1); -- 
    cr_3784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => type_cast_1231_inst_req_1); -- 
    cr_3676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => LOAD_out_depth_high_1203_load_0_req_1); -- 
    rr_3632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => LOAD_depth_high_1200_load_0_req_0); -- 
    cr_3770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => type_cast_1227_inst_req_1); -- 
    rr_3665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => LOAD_out_depth_high_1203_load_0_req_0); -- 
    cr_3709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => LOAD_out_col_high_1206_load_0_req_1); -- 
    cr_3610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => LOAD_pad_1197_load_0_req_1); -- 
    cr_3742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => type_cast_1214_inst_req_1); -- 
    rr_3599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => LOAD_pad_1197_load_0_req_0); -- 
    rr_3698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => LOAD_out_col_high_1206_load_0_req_0); -- 
    cr_3756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => type_cast_1218_inst_req_1); -- 
    cr_3728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => type_cast_1210_inst_req_1); -- 
    cr_3582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => type_cast_1188_inst_req_1); -- 
    rr_3577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(850), ack => type_cast_1188_inst_req_0); -- 
    zeropad3D_cp_element_group_850: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_850"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(848) & zeropad3D_CP_2067_elements(849);
      gj_zeropad3D_cp_element_group_850 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(850), clk => clk, reset => reset); --
    end block;
    -- CP-element group 851:  transition  input  bypass 
    -- CP-element group 851: predecessors 
    -- CP-element group 851: 	2 
    -- CP-element group 851: successors 
    -- CP-element group 851: 	853 
    -- CP-element group 851:  members (2) 
      -- CP-element group 851: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/Sample/$exit
      -- CP-element group 851: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/Sample/ra
      -- 
    ra_11070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 851_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1281_inst_ack_0, ack => zeropad3D_CP_2067_elements(851)); -- 
    -- CP-element group 852:  transition  input  bypass 
    -- CP-element group 852: predecessors 
    -- CP-element group 852: 	2 
    -- CP-element group 852: successors 
    -- CP-element group 852: 	853 
    -- CP-element group 852:  members (2) 
      -- CP-element group 852: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/Update/$exit
      -- CP-element group 852: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/Update/ca
      -- 
    ca_11075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 852_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1281_inst_ack_1, ack => zeropad3D_CP_2067_elements(852)); -- 
    -- CP-element group 853:  join  transition  output  bypass 
    -- CP-element group 853: predecessors 
    -- CP-element group 853: 	851 
    -- CP-element group 853: 	852 
    -- CP-element group 853: successors 
    -- CP-element group 853: 	860 
    -- CP-element group 853:  members (5) 
      -- CP-element group 853: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/$exit
      -- CP-element group 853: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/$exit
      -- CP-element group 853: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/$exit
      -- CP-element group 853: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1281/SplitProtocol/$exit
      -- CP-element group 853: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_req
      -- 
    phi_stmt_1276_req_11076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1276_req_11076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(853), ack => phi_stmt_1276_req_1); -- 
    zeropad3D_cp_element_group_853: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_853"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(851) & zeropad3D_CP_2067_elements(852);
      gj_zeropad3D_cp_element_group_853 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(853), clk => clk, reset => reset); --
    end block;
    -- CP-element group 854:  transition  input  bypass 
    -- CP-element group 854: predecessors 
    -- CP-element group 854: 	2 
    -- CP-element group 854: successors 
    -- CP-element group 854: 	856 
    -- CP-element group 854:  members (2) 
      -- CP-element group 854: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/Sample/$exit
      -- CP-element group 854: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/Sample/ra
      -- 
    ra_11093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 854_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1288_inst_ack_0, ack => zeropad3D_CP_2067_elements(854)); -- 
    -- CP-element group 855:  transition  input  bypass 
    -- CP-element group 855: predecessors 
    -- CP-element group 855: 	2 
    -- CP-element group 855: successors 
    -- CP-element group 855: 	856 
    -- CP-element group 855:  members (2) 
      -- CP-element group 855: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/Update/$exit
      -- CP-element group 855: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/Update/ca
      -- 
    ca_11098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 855_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1288_inst_ack_1, ack => zeropad3D_CP_2067_elements(855)); -- 
    -- CP-element group 856:  join  transition  output  bypass 
    -- CP-element group 856: predecessors 
    -- CP-element group 856: 	854 
    -- CP-element group 856: 	855 
    -- CP-element group 856: successors 
    -- CP-element group 856: 	860 
    -- CP-element group 856:  members (5) 
      -- CP-element group 856: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/$exit
      -- CP-element group 856: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/$exit
      -- CP-element group 856: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/$exit
      -- CP-element group 856: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1288/SplitProtocol/$exit
      -- CP-element group 856: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_req
      -- 
    phi_stmt_1282_req_11099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1282_req_11099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(856), ack => phi_stmt_1282_req_1); -- 
    zeropad3D_cp_element_group_856: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_856"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(854) & zeropad3D_CP_2067_elements(855);
      gj_zeropad3D_cp_element_group_856 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(856), clk => clk, reset => reset); --
    end block;
    -- CP-element group 857:  transition  input  bypass 
    -- CP-element group 857: predecessors 
    -- CP-element group 857: 	2 
    -- CP-element group 857: successors 
    -- CP-element group 857: 	859 
    -- CP-element group 857:  members (2) 
      -- CP-element group 857: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Sample/$exit
      -- CP-element group 857: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Sample/ra
      -- 
    ra_11116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 857_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1295_inst_ack_0, ack => zeropad3D_CP_2067_elements(857)); -- 
    -- CP-element group 858:  transition  input  bypass 
    -- CP-element group 858: predecessors 
    -- CP-element group 858: 	2 
    -- CP-element group 858: successors 
    -- CP-element group 858: 	859 
    -- CP-element group 858:  members (2) 
      -- CP-element group 858: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Update/$exit
      -- CP-element group 858: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Update/ca
      -- 
    ca_11121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 858_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1295_inst_ack_1, ack => zeropad3D_CP_2067_elements(858)); -- 
    -- CP-element group 859:  join  transition  output  bypass 
    -- CP-element group 859: predecessors 
    -- CP-element group 859: 	857 
    -- CP-element group 859: 	858 
    -- CP-element group 859: successors 
    -- CP-element group 859: 	860 
    -- CP-element group 859:  members (5) 
      -- CP-element group 859: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/$exit
      -- CP-element group 859: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/$exit
      -- CP-element group 859: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/$exit
      -- CP-element group 859: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/$exit
      -- CP-element group 859: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_req
      -- 
    phi_stmt_1289_req_11122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1289_req_11122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(859), ack => phi_stmt_1289_req_1); -- 
    zeropad3D_cp_element_group_859: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_859"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(857) & zeropad3D_CP_2067_elements(858);
      gj_zeropad3D_cp_element_group_859 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(859), clk => clk, reset => reset); --
    end block;
    -- CP-element group 860:  join  transition  bypass 
    -- CP-element group 860: predecessors 
    -- CP-element group 860: 	853 
    -- CP-element group 860: 	856 
    -- CP-element group 860: 	859 
    -- CP-element group 860: successors 
    -- CP-element group 860: 	867 
    -- CP-element group 860:  members (1) 
      -- CP-element group 860: 	 branch_block_stmt_655/ifx_xend389_whilex_xbody234_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_860: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_860"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(853) & zeropad3D_CP_2067_elements(856) & zeropad3D_CP_2067_elements(859);
      gj_zeropad3D_cp_element_group_860 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(860), clk => clk, reset => reset); --
    end block;
    -- CP-element group 861:  transition  input  bypass 
    -- CP-element group 861: predecessors 
    -- CP-element group 861: 	130 
    -- CP-element group 861: successors 
    -- CP-element group 861: 	863 
    -- CP-element group 861:  members (2) 
      -- CP-element group 861: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/Sample/$exit
      -- CP-element group 861: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/Sample/ra
      -- 
    ra_11142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 861_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_0, ack => zeropad3D_CP_2067_elements(861)); -- 
    -- CP-element group 862:  transition  input  bypass 
    -- CP-element group 862: predecessors 
    -- CP-element group 862: 	130 
    -- CP-element group 862: successors 
    -- CP-element group 862: 	863 
    -- CP-element group 862:  members (2) 
      -- CP-element group 862: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/Update/$exit
      -- CP-element group 862: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/Update/ca
      -- 
    ca_11147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 862_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_1, ack => zeropad3D_CP_2067_elements(862)); -- 
    -- CP-element group 863:  join  transition  output  bypass 
    -- CP-element group 863: predecessors 
    -- CP-element group 863: 	861 
    -- CP-element group 863: 	862 
    -- CP-element group 863: successors 
    -- CP-element group 863: 	866 
    -- CP-element group 863:  members (5) 
      -- CP-element group 863: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/$exit
      -- CP-element group 863: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/$exit
      -- CP-element group 863: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/$exit
      -- CP-element group 863: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_sources/type_cast_1279/SplitProtocol/$exit
      -- CP-element group 863: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1276/phi_stmt_1276_req
      -- 
    phi_stmt_1276_req_11148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1276_req_11148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(863), ack => phi_stmt_1276_req_0); -- 
    zeropad3D_cp_element_group_863: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_863"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(861) & zeropad3D_CP_2067_elements(862);
      gj_zeropad3D_cp_element_group_863 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(863), clk => clk, reset => reset); --
    end block;
    -- CP-element group 864:  transition  output  delay-element  bypass 
    -- CP-element group 864: predecessors 
    -- CP-element group 864: 	130 
    -- CP-element group 864: successors 
    -- CP-element group 864: 	866 
    -- CP-element group 864:  members (4) 
      -- CP-element group 864: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1282/$exit
      -- CP-element group 864: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/$exit
      -- CP-element group 864: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_sources/type_cast_1286_konst_delay_trans
      -- CP-element group 864: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1282/phi_stmt_1282_req
      -- 
    phi_stmt_1282_req_11156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1282_req_11156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(864), ack => phi_stmt_1282_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(864) is a control-delay.
    cp_element_864_delay: control_delay_element  generic map(name => " 864_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(130), ack => zeropad3D_CP_2067_elements(864), clk => clk, reset =>reset);
    -- CP-element group 865:  transition  output  delay-element  bypass 
    -- CP-element group 865: predecessors 
    -- CP-element group 865: 	130 
    -- CP-element group 865: successors 
    -- CP-element group 865: 	866 
    -- CP-element group 865:  members (4) 
      -- CP-element group 865: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1289/$exit
      -- CP-element group 865: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/$exit
      -- CP-element group 865: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1293_konst_delay_trans
      -- CP-element group 865: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/phi_stmt_1289/phi_stmt_1289_req
      -- 
    phi_stmt_1289_req_11164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1289_req_11164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(865), ack => phi_stmt_1289_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(865) is a control-delay.
    cp_element_865_delay: control_delay_element  generic map(name => " 865_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(130), ack => zeropad3D_CP_2067_elements(865), clk => clk, reset =>reset);
    -- CP-element group 866:  join  transition  bypass 
    -- CP-element group 866: predecessors 
    -- CP-element group 866: 	863 
    -- CP-element group 866: 	864 
    -- CP-element group 866: 	865 
    -- CP-element group 866: successors 
    -- CP-element group 866: 	867 
    -- CP-element group 866:  members (1) 
      -- CP-element group 866: 	 branch_block_stmt_655/whilex_xend_whilex_xbody234_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_866: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_866"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(863) & zeropad3D_CP_2067_elements(864) & zeropad3D_CP_2067_elements(865);
      gj_zeropad3D_cp_element_group_866 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(866), clk => clk, reset => reset); --
    end block;
    -- CP-element group 867:  merge  fork  transition  place  bypass 
    -- CP-element group 867: predecessors 
    -- CP-element group 867: 	860 
    -- CP-element group 867: 	866 
    -- CP-element group 867: successors 
    -- CP-element group 867: 	868 
    -- CP-element group 867: 	869 
    -- CP-element group 867: 	870 
    -- CP-element group 867:  members (2) 
      -- CP-element group 867: 	 branch_block_stmt_655/merge_stmt_1275_PhiReqMerge
      -- CP-element group 867: 	 branch_block_stmt_655/merge_stmt_1275_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(867) <= OrReduce(zeropad3D_CP_2067_elements(860) & zeropad3D_CP_2067_elements(866));
    -- CP-element group 868:  transition  input  bypass 
    -- CP-element group 868: predecessors 
    -- CP-element group 868: 	867 
    -- CP-element group 868: successors 
    -- CP-element group 868: 	871 
    -- CP-element group 868:  members (1) 
      -- CP-element group 868: 	 branch_block_stmt_655/merge_stmt_1275_PhiAck/phi_stmt_1276_ack
      -- 
    phi_stmt_1276_ack_11169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 868_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1276_ack_0, ack => zeropad3D_CP_2067_elements(868)); -- 
    -- CP-element group 869:  transition  input  bypass 
    -- CP-element group 869: predecessors 
    -- CP-element group 869: 	867 
    -- CP-element group 869: successors 
    -- CP-element group 869: 	871 
    -- CP-element group 869:  members (1) 
      -- CP-element group 869: 	 branch_block_stmt_655/merge_stmt_1275_PhiAck/phi_stmt_1282_ack
      -- 
    phi_stmt_1282_ack_11170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 869_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1282_ack_0, ack => zeropad3D_CP_2067_elements(869)); -- 
    -- CP-element group 870:  transition  input  bypass 
    -- CP-element group 870: predecessors 
    -- CP-element group 870: 	867 
    -- CP-element group 870: successors 
    -- CP-element group 870: 	871 
    -- CP-element group 870:  members (1) 
      -- CP-element group 870: 	 branch_block_stmt_655/merge_stmt_1275_PhiAck/phi_stmt_1289_ack
      -- 
    phi_stmt_1289_ack_11171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 870_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1289_ack_0, ack => zeropad3D_CP_2067_elements(870)); -- 
    -- CP-element group 871:  join  fork  transition  place  output  bypass 
    -- CP-element group 871: predecessors 
    -- CP-element group 871: 	868 
    -- CP-element group 871: 	869 
    -- CP-element group 871: 	870 
    -- CP-element group 871: successors 
    -- CP-element group 871: 	131 
    -- CP-element group 871: 	132 
    -- CP-element group 871:  members (10) 
      -- CP-element group 871: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_Sample/rr
      -- CP-element group 871: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/$entry
      -- CP-element group 871: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_Update/$entry
      -- CP-element group 871: 	 branch_block_stmt_655/merge_stmt_1275__exit__
      -- CP-element group 871: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308__entry__
      -- CP-element group 871: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_Update/cr
      -- CP-element group 871: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_Sample/$entry
      -- CP-element group 871: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_update_start_
      -- CP-element group 871: 	 branch_block_stmt_655/assign_stmt_1301_to_assign_stmt_1308/type_cast_1300_sample_start_
      -- CP-element group 871: 	 branch_block_stmt_655/merge_stmt_1275_PhiAck/$exit
      -- 
    rr_3796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(871), ack => type_cast_1300_inst_req_0); -- 
    cr_3801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(871), ack => type_cast_1300_inst_req_1); -- 
    zeropad3D_cp_element_group_871: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_871"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(868) & zeropad3D_CP_2067_elements(869) & zeropad3D_CP_2067_elements(870);
      gj_zeropad3D_cp_element_group_871 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(871), clk => clk, reset => reset); --
    end block;
    -- CP-element group 872:  merge  fork  transition  place  output  bypass 
    -- CP-element group 872: predecessors 
    -- CP-element group 872: 	133 
    -- CP-element group 872: 	140 
    -- CP-element group 872: 	143 
    -- CP-element group 872: 	150 
    -- CP-element group 872: successors 
    -- CP-element group 872: 	151 
    -- CP-element group 872: 	152 
    -- CP-element group 872: 	153 
    -- CP-element group 872: 	154 
    -- CP-element group 872: 	157 
    -- CP-element group 872: 	159 
    -- CP-element group 872: 	161 
    -- CP-element group 872: 	163 
    -- CP-element group 872:  members (33) 
      -- CP-element group 872: 	 branch_block_stmt_655/merge_stmt_1392__exit__
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448__entry__
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_sample_start_
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_update_start_
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_Sample/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_Sample/rr
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_Update/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1396_Update/cr
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_sample_start_
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_update_start_
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_Sample/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_Sample/rr
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_Update/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1401_Update/cr
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_update_start_
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_Update/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/type_cast_1435_Update/cr
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_update_start_
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_update_start
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_Update/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/array_obj_ref_1441_final_index_sum_regn_Update/req
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_complete/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/addr_of_1442_complete/req
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_update_start_
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Update/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Update/word_access_complete/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Update/word_access_complete/word_0/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/assign_stmt_1397_to_assign_stmt_1448/ptr_deref_1445_Update/word_access_complete/word_0/cr
      -- CP-element group 872: 	 branch_block_stmt_655/merge_stmt_1392_PhiReqMerge
      -- CP-element group 872: 	 branch_block_stmt_655/merge_stmt_1392_PhiAck/$entry
      -- CP-element group 872: 	 branch_block_stmt_655/merge_stmt_1392_PhiAck/$exit
      -- CP-element group 872: 	 branch_block_stmt_655/merge_stmt_1392_PhiAck/dummy
      -- 
    rr_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(872), ack => type_cast_1396_inst_req_0); -- 
    cr_4011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(872), ack => type_cast_1396_inst_req_1); -- 
    rr_4020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(872), ack => type_cast_1401_inst_req_0); -- 
    cr_4025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(872), ack => type_cast_1401_inst_req_1); -- 
    cr_4039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(872), ack => type_cast_1435_inst_req_1); -- 
    req_4070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(872), ack => array_obj_ref_1441_index_offset_req_1); -- 
    req_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(872), ack => addr_of_1442_final_reg_req_1); -- 
    cr_4135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(872), ack => ptr_deref_1445_store_0_req_1); -- 
    zeropad3D_CP_2067_elements(872) <= OrReduce(zeropad3D_CP_2067_elements(133) & zeropad3D_CP_2067_elements(140) & zeropad3D_CP_2067_elements(143) & zeropad3D_CP_2067_elements(150));
    -- CP-element group 873:  merge  fork  transition  place  output  bypass 
    -- CP-element group 873: predecessors 
    -- CP-element group 873: 	164 
    -- CP-element group 873: 	184 
    -- CP-element group 873: successors 
    -- CP-element group 873: 	185 
    -- CP-element group 873: 	186 
    -- CP-element group 873:  members (13) 
      -- CP-element group 873: 	 branch_block_stmt_655/merge_stmt_1557__exit__
      -- CP-element group 873: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575__entry__
      -- CP-element group 873: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/$entry
      -- CP-element group 873: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_sample_start_
      -- CP-element group 873: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_update_start_
      -- CP-element group 873: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_Sample/$entry
      -- CP-element group 873: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_Sample/rr
      -- CP-element group 873: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_Update/$entry
      -- CP-element group 873: 	 branch_block_stmt_655/assign_stmt_1562_to_assign_stmt_1575/type_cast_1561_Update/cr
      -- CP-element group 873: 	 branch_block_stmt_655/merge_stmt_1557_PhiAck/dummy
      -- CP-element group 873: 	 branch_block_stmt_655/merge_stmt_1557_PhiAck/$exit
      -- CP-element group 873: 	 branch_block_stmt_655/merge_stmt_1557_PhiAck/$entry
      -- CP-element group 873: 	 branch_block_stmt_655/merge_stmt_1557_PhiReqMerge
      -- 
    rr_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(873), ack => type_cast_1561_inst_req_0); -- 
    cr_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(873), ack => type_cast_1561_inst_req_1); -- 
    zeropad3D_CP_2067_elements(873) <= OrReduce(zeropad3D_CP_2067_elements(164) & zeropad3D_CP_2067_elements(184));
    -- CP-element group 874:  transition  output  delay-element  bypass 
    -- CP-element group 874: predecessors 
    -- CP-element group 874: 	206 
    -- CP-element group 874: successors 
    -- CP-element group 874: 	881 
    -- CP-element group 874:  members (4) 
      -- CP-element group 874: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_req
      -- CP-element group 874: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1687_konst_delay_trans
      -- CP-element group 874: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/$exit
      -- CP-element group 874: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1681/$exit
      -- 
    phi_stmt_1681_req_11282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1681_req_11282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(874), ack => phi_stmt_1681_req_1); -- 
    -- Element group zeropad3D_CP_2067_elements(874) is a control-delay.
    cp_element_874_delay: control_delay_element  generic map(name => " 874_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(206), ack => zeropad3D_CP_2067_elements(874), clk => clk, reset =>reset);
    -- CP-element group 875:  transition  input  bypass 
    -- CP-element group 875: predecessors 
    -- CP-element group 875: 	206 
    -- CP-element group 875: successors 
    -- CP-element group 875: 	877 
    -- CP-element group 875:  members (2) 
      -- CP-element group 875: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/Sample/ra
      -- CP-element group 875: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/Sample/$exit
      -- 
    ra_11299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 875_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1678_inst_ack_0, ack => zeropad3D_CP_2067_elements(875)); -- 
    -- CP-element group 876:  transition  input  bypass 
    -- CP-element group 876: predecessors 
    -- CP-element group 876: 	206 
    -- CP-element group 876: successors 
    -- CP-element group 876: 	877 
    -- CP-element group 876:  members (2) 
      -- CP-element group 876: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/Update/ca
      -- CP-element group 876: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/Update/$exit
      -- 
    ca_11304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 876_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1678_inst_ack_1, ack => zeropad3D_CP_2067_elements(876)); -- 
    -- CP-element group 877:  join  transition  output  bypass 
    -- CP-element group 877: predecessors 
    -- CP-element group 877: 	875 
    -- CP-element group 877: 	876 
    -- CP-element group 877: successors 
    -- CP-element group 877: 	881 
    -- CP-element group 877:  members (5) 
      -- CP-element group 877: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/$exit
      -- CP-element group 877: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1678/SplitProtocol/$exit
      -- CP-element group 877: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/$exit
      -- CP-element group 877: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/$exit
      -- CP-element group 877: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_req
      -- 
    phi_stmt_1675_req_11305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1675_req_11305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(877), ack => phi_stmt_1675_req_0); -- 
    zeropad3D_cp_element_group_877: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_877"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(875) & zeropad3D_CP_2067_elements(876);
      gj_zeropad3D_cp_element_group_877 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(877), clk => clk, reset => reset); --
    end block;
    -- CP-element group 878:  transition  input  bypass 
    -- CP-element group 878: predecessors 
    -- CP-element group 878: 	206 
    -- CP-element group 878: successors 
    -- CP-element group 878: 	880 
    -- CP-element group 878:  members (2) 
      -- CP-element group 878: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/Sample/$exit
      -- CP-element group 878: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/Sample/ra
      -- 
    ra_11322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 878_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1674_inst_ack_0, ack => zeropad3D_CP_2067_elements(878)); -- 
    -- CP-element group 879:  transition  input  bypass 
    -- CP-element group 879: predecessors 
    -- CP-element group 879: 	206 
    -- CP-element group 879: successors 
    -- CP-element group 879: 	880 
    -- CP-element group 879:  members (2) 
      -- CP-element group 879: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/Update/ca
      -- CP-element group 879: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/Update/$exit
      -- 
    ca_11327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 879_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1674_inst_ack_1, ack => zeropad3D_CP_2067_elements(879)); -- 
    -- CP-element group 880:  join  transition  output  bypass 
    -- CP-element group 880: predecessors 
    -- CP-element group 880: 	878 
    -- CP-element group 880: 	879 
    -- CP-element group 880: successors 
    -- CP-element group 880: 	881 
    -- CP-element group 880:  members (5) 
      -- CP-element group 880: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_req
      -- CP-element group 880: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/$exit
      -- CP-element group 880: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/$exit
      -- CP-element group 880: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/$exit
      -- CP-element group 880: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1674/SplitProtocol/$exit
      -- 
    phi_stmt_1669_req_11328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1669_req_11328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(880), ack => phi_stmt_1669_req_1); -- 
    zeropad3D_cp_element_group_880: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_880"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(878) & zeropad3D_CP_2067_elements(879);
      gj_zeropad3D_cp_element_group_880 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(880), clk => clk, reset => reset); --
    end block;
    -- CP-element group 881:  join  transition  bypass 
    -- CP-element group 881: predecessors 
    -- CP-element group 881: 	874 
    -- CP-element group 881: 	877 
    -- CP-element group 881: 	880 
    -- CP-element group 881: successors 
    -- CP-element group 881: 	892 
    -- CP-element group 881:  members (1) 
      -- CP-element group 881: 	 branch_block_stmt_655/ifx_xelse353_ifx_xend389_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_881: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_881"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(874) & zeropad3D_CP_2067_elements(877) & zeropad3D_CP_2067_elements(880);
      gj_zeropad3D_cp_element_group_881 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(881), clk => clk, reset => reset); --
    end block;
    -- CP-element group 882:  transition  input  bypass 
    -- CP-element group 882: predecessors 
    -- CP-element group 882: 	187 
    -- CP-element group 882: successors 
    -- CP-element group 882: 	884 
    -- CP-element group 882:  members (2) 
      -- CP-element group 882: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/Sample/ra
      -- CP-element group 882: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/Sample/$exit
      -- 
    ra_11348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 882_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1684_inst_ack_0, ack => zeropad3D_CP_2067_elements(882)); -- 
    -- CP-element group 883:  transition  input  bypass 
    -- CP-element group 883: predecessors 
    -- CP-element group 883: 	187 
    -- CP-element group 883: successors 
    -- CP-element group 883: 	884 
    -- CP-element group 883:  members (2) 
      -- CP-element group 883: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/Update/ca
      -- CP-element group 883: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/Update/$exit
      -- 
    ca_11353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 883_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1684_inst_ack_1, ack => zeropad3D_CP_2067_elements(883)); -- 
    -- CP-element group 884:  join  transition  output  bypass 
    -- CP-element group 884: predecessors 
    -- CP-element group 884: 	882 
    -- CP-element group 884: 	883 
    -- CP-element group 884: successors 
    -- CP-element group 884: 	891 
    -- CP-element group 884:  members (5) 
      -- CP-element group 884: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_req
      -- CP-element group 884: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/SplitProtocol/$exit
      -- CP-element group 884: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/type_cast_1684/$exit
      -- CP-element group 884: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/phi_stmt_1681_sources/$exit
      -- CP-element group 884: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1681/$exit
      -- 
    phi_stmt_1681_req_11354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1681_req_11354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(884), ack => phi_stmt_1681_req_0); -- 
    zeropad3D_cp_element_group_884: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_884"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(882) & zeropad3D_CP_2067_elements(883);
      gj_zeropad3D_cp_element_group_884 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(884), clk => clk, reset => reset); --
    end block;
    -- CP-element group 885:  transition  input  bypass 
    -- CP-element group 885: predecessors 
    -- CP-element group 885: 	187 
    -- CP-element group 885: successors 
    -- CP-element group 885: 	887 
    -- CP-element group 885:  members (2) 
      -- CP-element group 885: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/Sample/$exit
      -- CP-element group 885: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/Sample/ra
      -- 
    ra_11371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 885_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1680_inst_ack_0, ack => zeropad3D_CP_2067_elements(885)); -- 
    -- CP-element group 886:  transition  input  bypass 
    -- CP-element group 886: predecessors 
    -- CP-element group 886: 	187 
    -- CP-element group 886: successors 
    -- CP-element group 886: 	887 
    -- CP-element group 886:  members (2) 
      -- CP-element group 886: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/Update/$exit
      -- CP-element group 886: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/Update/ca
      -- 
    ca_11376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 886_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1680_inst_ack_1, ack => zeropad3D_CP_2067_elements(886)); -- 
    -- CP-element group 887:  join  transition  output  bypass 
    -- CP-element group 887: predecessors 
    -- CP-element group 887: 	885 
    -- CP-element group 887: 	886 
    -- CP-element group 887: successors 
    -- CP-element group 887: 	891 
    -- CP-element group 887:  members (5) 
      -- CP-element group 887: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_req
      -- CP-element group 887: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/SplitProtocol/$exit
      -- CP-element group 887: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/type_cast_1680/$exit
      -- CP-element group 887: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/phi_stmt_1675_sources/$exit
      -- CP-element group 887: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1675/$exit
      -- 
    phi_stmt_1675_req_11377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1675_req_11377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(887), ack => phi_stmt_1675_req_1); -- 
    zeropad3D_cp_element_group_887: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_887"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(885) & zeropad3D_CP_2067_elements(886);
      gj_zeropad3D_cp_element_group_887 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(887), clk => clk, reset => reset); --
    end block;
    -- CP-element group 888:  transition  input  bypass 
    -- CP-element group 888: predecessors 
    -- CP-element group 888: 	187 
    -- CP-element group 888: successors 
    -- CP-element group 888: 	890 
    -- CP-element group 888:  members (2) 
      -- CP-element group 888: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/Sample/ra
      -- CP-element group 888: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/Sample/$exit
      -- 
    ra_11394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 888_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_0, ack => zeropad3D_CP_2067_elements(888)); -- 
    -- CP-element group 889:  transition  input  bypass 
    -- CP-element group 889: predecessors 
    -- CP-element group 889: 	187 
    -- CP-element group 889: successors 
    -- CP-element group 889: 	890 
    -- CP-element group 889:  members (2) 
      -- CP-element group 889: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/Update/ca
      -- CP-element group 889: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/Update/$exit
      -- 
    ca_11399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 889_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_1, ack => zeropad3D_CP_2067_elements(889)); -- 
    -- CP-element group 890:  join  transition  output  bypass 
    -- CP-element group 890: predecessors 
    -- CP-element group 890: 	888 
    -- CP-element group 890: 	889 
    -- CP-element group 890: successors 
    -- CP-element group 890: 	891 
    -- CP-element group 890:  members (5) 
      -- CP-element group 890: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/$exit
      -- CP-element group 890: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_req
      -- CP-element group 890: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/SplitProtocol/$exit
      -- CP-element group 890: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/type_cast_1672/$exit
      -- CP-element group 890: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/phi_stmt_1669/phi_stmt_1669_sources/$exit
      -- 
    phi_stmt_1669_req_11400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1669_req_11400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(890), ack => phi_stmt_1669_req_0); -- 
    zeropad3D_cp_element_group_890: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_890"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(888) & zeropad3D_CP_2067_elements(889);
      gj_zeropad3D_cp_element_group_890 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(890), clk => clk, reset => reset); --
    end block;
    -- CP-element group 891:  join  transition  bypass 
    -- CP-element group 891: predecessors 
    -- CP-element group 891: 	884 
    -- CP-element group 891: 	887 
    -- CP-element group 891: 	890 
    -- CP-element group 891: successors 
    -- CP-element group 891: 	892 
    -- CP-element group 891:  members (1) 
      -- CP-element group 891: 	 branch_block_stmt_655/ifx_xthen348_ifx_xend389_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_891: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_891"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(884) & zeropad3D_CP_2067_elements(887) & zeropad3D_CP_2067_elements(890);
      gj_zeropad3D_cp_element_group_891 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(891), clk => clk, reset => reset); --
    end block;
    -- CP-element group 892:  merge  fork  transition  place  bypass 
    -- CP-element group 892: predecessors 
    -- CP-element group 892: 	881 
    -- CP-element group 892: 	891 
    -- CP-element group 892: successors 
    -- CP-element group 892: 	893 
    -- CP-element group 892: 	894 
    -- CP-element group 892: 	895 
    -- CP-element group 892:  members (2) 
      -- CP-element group 892: 	 branch_block_stmt_655/merge_stmt_1668_PhiReqMerge
      -- CP-element group 892: 	 branch_block_stmt_655/merge_stmt_1668_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(892) <= OrReduce(zeropad3D_CP_2067_elements(881) & zeropad3D_CP_2067_elements(891));
    -- CP-element group 893:  transition  input  bypass 
    -- CP-element group 893: predecessors 
    -- CP-element group 893: 	892 
    -- CP-element group 893: successors 
    -- CP-element group 893: 	896 
    -- CP-element group 893:  members (1) 
      -- CP-element group 893: 	 branch_block_stmt_655/merge_stmt_1668_PhiAck/phi_stmt_1669_ack
      -- 
    phi_stmt_1669_ack_11405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 893_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1669_ack_0, ack => zeropad3D_CP_2067_elements(893)); -- 
    -- CP-element group 894:  transition  input  bypass 
    -- CP-element group 894: predecessors 
    -- CP-element group 894: 	892 
    -- CP-element group 894: successors 
    -- CP-element group 894: 	896 
    -- CP-element group 894:  members (1) 
      -- CP-element group 894: 	 branch_block_stmt_655/merge_stmt_1668_PhiAck/phi_stmt_1675_ack
      -- 
    phi_stmt_1675_ack_11406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 894_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1675_ack_0, ack => zeropad3D_CP_2067_elements(894)); -- 
    -- CP-element group 895:  transition  input  bypass 
    -- CP-element group 895: predecessors 
    -- CP-element group 895: 	892 
    -- CP-element group 895: successors 
    -- CP-element group 895: 	896 
    -- CP-element group 895:  members (1) 
      -- CP-element group 895: 	 branch_block_stmt_655/merge_stmt_1668_PhiAck/phi_stmt_1681_ack
      -- 
    phi_stmt_1681_ack_11407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 895_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1681_ack_0, ack => zeropad3D_CP_2067_elements(895)); -- 
    -- CP-element group 896:  join  transition  bypass 
    -- CP-element group 896: predecessors 
    -- CP-element group 896: 	893 
    -- CP-element group 896: 	894 
    -- CP-element group 896: 	895 
    -- CP-element group 896: successors 
    -- CP-element group 896: 	2 
    -- CP-element group 896:  members (1) 
      -- CP-element group 896: 	 branch_block_stmt_655/merge_stmt_1668_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_896: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_896"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(893) & zeropad3D_CP_2067_elements(894) & zeropad3D_CP_2067_elements(895);
      gj_zeropad3D_cp_element_group_896 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(896), clk => clk, reset => reset); --
    end block;
    -- CP-element group 897:  transition  input  bypass 
    -- CP-element group 897: predecessors 
    -- CP-element group 897: 	205 
    -- CP-element group 897: successors 
    -- CP-element group 897: 	899 
    -- CP-element group 897:  members (2) 
      -- CP-element group 897: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/Sample/ra
      -- CP-element group 897: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/Sample/$exit
      -- 
    ra_11427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 897_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1698_inst_ack_0, ack => zeropad3D_CP_2067_elements(897)); -- 
    -- CP-element group 898:  transition  input  bypass 
    -- CP-element group 898: predecessors 
    -- CP-element group 898: 	205 
    -- CP-element group 898: successors 
    -- CP-element group 898: 	899 
    -- CP-element group 898:  members (2) 
      -- CP-element group 898: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/Update/ca
      -- CP-element group 898: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/Update/$exit
      -- 
    ca_11432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 898_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1698_inst_ack_1, ack => zeropad3D_CP_2067_elements(898)); -- 
    -- CP-element group 899:  join  transition  output  bypass 
    -- CP-element group 899: predecessors 
    -- CP-element group 899: 	897 
    -- CP-element group 899: 	898 
    -- CP-element group 899: successors 
    -- CP-element group 899: 	903 
    -- CP-element group 899:  members (5) 
      -- CP-element group 899: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/$exit
      -- CP-element group 899: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_req
      -- CP-element group 899: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/SplitProtocol/$exit
      -- CP-element group 899: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/type_cast_1698/$exit
      -- CP-element group 899: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1695/phi_stmt_1695_sources/$exit
      -- 
    phi_stmt_1695_req_11433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1695_req_11433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(899), ack => phi_stmt_1695_req_0); -- 
    zeropad3D_cp_element_group_899: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_899"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(897) & zeropad3D_CP_2067_elements(898);
      gj_zeropad3D_cp_element_group_899 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(899), clk => clk, reset => reset); --
    end block;
    -- CP-element group 900:  transition  input  bypass 
    -- CP-element group 900: predecessors 
    -- CP-element group 900: 	205 
    -- CP-element group 900: successors 
    -- CP-element group 900: 	902 
    -- CP-element group 900:  members (2) 
      -- CP-element group 900: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/Sample/ra
      -- CP-element group 900: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/Sample/$exit
      -- 
    ra_11450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 900_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1694_inst_ack_0, ack => zeropad3D_CP_2067_elements(900)); -- 
    -- CP-element group 901:  transition  input  bypass 
    -- CP-element group 901: predecessors 
    -- CP-element group 901: 	205 
    -- CP-element group 901: successors 
    -- CP-element group 901: 	902 
    -- CP-element group 901:  members (2) 
      -- CP-element group 901: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/Update/ca
      -- CP-element group 901: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/Update/$exit
      -- 
    ca_11455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 901_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1694_inst_ack_1, ack => zeropad3D_CP_2067_elements(901)); -- 
    -- CP-element group 902:  join  transition  output  bypass 
    -- CP-element group 902: predecessors 
    -- CP-element group 902: 	900 
    -- CP-element group 902: 	901 
    -- CP-element group 902: successors 
    -- CP-element group 902: 	903 
    -- CP-element group 902:  members (5) 
      -- CP-element group 902: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_req
      -- CP-element group 902: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/SplitProtocol/$exit
      -- CP-element group 902: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/type_cast_1694/$exit
      -- CP-element group 902: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/phi_stmt_1691_sources/$exit
      -- CP-element group 902: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/phi_stmt_1691/$exit
      -- 
    phi_stmt_1691_req_11456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1691_req_11456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(902), ack => phi_stmt_1691_req_0); -- 
    zeropad3D_cp_element_group_902: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_902"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(900) & zeropad3D_CP_2067_elements(901);
      gj_zeropad3D_cp_element_group_902 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(902), clk => clk, reset => reset); --
    end block;
    -- CP-element group 903:  join  fork  transition  place  bypass 
    -- CP-element group 903: predecessors 
    -- CP-element group 903: 	899 
    -- CP-element group 903: 	902 
    -- CP-element group 903: successors 
    -- CP-element group 903: 	904 
    -- CP-element group 903: 	905 
    -- CP-element group 903:  members (3) 
      -- CP-element group 903: 	 branch_block_stmt_655/merge_stmt_1690_PhiReqMerge
      -- CP-element group 903: 	 branch_block_stmt_655/ifx_xelse353_whilex_xend390_PhiReq/$exit
      -- CP-element group 903: 	 branch_block_stmt_655/merge_stmt_1690_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_903: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_903"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(899) & zeropad3D_CP_2067_elements(902);
      gj_zeropad3D_cp_element_group_903 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(903), clk => clk, reset => reset); --
    end block;
    -- CP-element group 904:  transition  input  bypass 
    -- CP-element group 904: predecessors 
    -- CP-element group 904: 	903 
    -- CP-element group 904: successors 
    -- CP-element group 904: 	906 
    -- CP-element group 904:  members (1) 
      -- CP-element group 904: 	 branch_block_stmt_655/merge_stmt_1690_PhiAck/phi_stmt_1691_ack
      -- 
    phi_stmt_1691_ack_11461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 904_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1691_ack_0, ack => zeropad3D_CP_2067_elements(904)); -- 
    -- CP-element group 905:  transition  input  bypass 
    -- CP-element group 905: predecessors 
    -- CP-element group 905: 	903 
    -- CP-element group 905: successors 
    -- CP-element group 905: 	906 
    -- CP-element group 905:  members (1) 
      -- CP-element group 905: 	 branch_block_stmt_655/merge_stmt_1690_PhiAck/phi_stmt_1695_ack
      -- 
    phi_stmt_1695_ack_11462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 905_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1695_ack_0, ack => zeropad3D_CP_2067_elements(905)); -- 
    -- CP-element group 906:  join  fork  transition  place  output  bypass 
    -- CP-element group 906: predecessors 
    -- CP-element group 906: 	904 
    -- CP-element group 906: 	905 
    -- CP-element group 906: successors 
    -- CP-element group 906: 	207 
    -- CP-element group 906: 	208 
    -- CP-element group 906: 	209 
    -- CP-element group 906: 	210 
    -- CP-element group 906: 	211 
    -- CP-element group 906: 	212 
    -- CP-element group 906: 	213 
    -- CP-element group 906: 	214 
    -- CP-element group 906: 	215 
    -- CP-element group 906: 	216 
    -- CP-element group 906: 	218 
    -- CP-element group 906: 	220 
    -- CP-element group 906: 	222 
    -- CP-element group 906: 	224 
    -- CP-element group 906: 	226 
    -- CP-element group 906:  members (73) 
      -- CP-element group 906: 	 branch_block_stmt_655/merge_stmt_1690__exit__
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787__entry__
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Sample/word_access_start/word_0/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_word_address_calculated
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_root_address_calculated
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Sample/word_access_start/word_0/rr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Sample/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/word_access_complete/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_Update/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Sample/word_access_start/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Sample/word_access_start/word_0/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/word_access_complete/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Sample/word_access_start/word_0/rr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/word_access_complete/word_0/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Sample/word_access_start/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Sample/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1732_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_root_address_calculated
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_word_address_calculated
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_Update/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_sample_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_sample_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1728_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_Update/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_Update/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_col_high_1720_Update/word_access_complete/word_0/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1745_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1724_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1741_Update/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/word_access_complete/word_0/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_out_depth_high_1717_Update/word_access_complete/word_0/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_sample_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_Sample/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_Sample/rr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/type_cast_1702_Update/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_sample_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_word_address_calculated
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_root_address_calculated
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Sample/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Sample/word_access_start/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Sample/word_access_start/word_0/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Sample/word_access_start/word_0/rr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/word_access_complete/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/word_access_complete/word_0/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_pad_1711_Update/word_access_complete/word_0/cr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_sample_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_update_start_
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_word_address_calculated
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_root_address_calculated
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Sample/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Sample/word_access_start/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Sample/word_access_start/word_0/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Sample/word_access_start/word_0/rr
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/word_access_complete/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/word_access_complete/word_0/$entry
      -- CP-element group 906: 	 branch_block_stmt_655/assign_stmt_1703_to_assign_stmt_1787/LOAD_depth_high_1714_Update/word_access_complete/word_0/cr
      -- CP-element group 906: 	 branch_block_stmt_655/merge_stmt_1690_PhiAck/$exit
      -- 
    rr_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => LOAD_out_col_high_1720_load_0_req_0); -- 
    cr_4760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => type_cast_1732_inst_req_1); -- 
    rr_4669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => LOAD_out_depth_high_1717_load_0_req_0); -- 
    cr_4746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => type_cast_1728_inst_req_1); -- 
    cr_4732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => type_cast_1724_inst_req_1); -- 
    cr_4788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => type_cast_1745_inst_req_1); -- 
    cr_4713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => LOAD_out_col_high_1720_load_0_req_1); -- 
    cr_4774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => type_cast_1741_inst_req_1); -- 
    cr_4680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => LOAD_out_depth_high_1717_load_0_req_1); -- 
    rr_4581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => type_cast_1702_inst_req_0); -- 
    cr_4586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => type_cast_1702_inst_req_1); -- 
    rr_4603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => LOAD_pad_1711_load_0_req_0); -- 
    cr_4614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => LOAD_pad_1711_load_0_req_1); -- 
    rr_4636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => LOAD_depth_high_1714_load_0_req_0); -- 
    cr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(906), ack => LOAD_depth_high_1714_load_0_req_1); -- 
    zeropad3D_cp_element_group_906: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_906"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(904) & zeropad3D_CP_2067_elements(905);
      gj_zeropad3D_cp_element_group_906 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(906), clk => clk, reset => reset); --
    end block;
    -- CP-element group 907:  transition  input  bypass 
    -- CP-element group 907: predecessors 
    -- CP-element group 907: 	3 
    -- CP-element group 907: successors 
    -- CP-element group 907: 	909 
    -- CP-element group 907:  members (2) 
      -- CP-element group 907: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Sample/$exit
      -- CP-element group 907: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Sample/ra
      -- 
    ra_11482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 907_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1809_inst_ack_0, ack => zeropad3D_CP_2067_elements(907)); -- 
    -- CP-element group 908:  transition  input  bypass 
    -- CP-element group 908: predecessors 
    -- CP-element group 908: 	3 
    -- CP-element group 908: successors 
    -- CP-element group 908: 	909 
    -- CP-element group 908:  members (2) 
      -- CP-element group 908: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Update/ca
      -- CP-element group 908: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Update/$exit
      -- 
    ca_11487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 908_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1809_inst_ack_1, ack => zeropad3D_CP_2067_elements(908)); -- 
    -- CP-element group 909:  join  transition  output  bypass 
    -- CP-element group 909: predecessors 
    -- CP-element group 909: 	907 
    -- CP-element group 909: 	908 
    -- CP-element group 909: successors 
    -- CP-element group 909: 	916 
    -- CP-element group 909:  members (5) 
      -- CP-element group 909: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/$exit
      -- CP-element group 909: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/$exit
      -- CP-element group 909: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$exit
      -- CP-element group 909: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/$exit
      -- CP-element group 909: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_req
      -- 
    phi_stmt_1803_req_11488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1803_req_11488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(909), ack => phi_stmt_1803_req_1); -- 
    zeropad3D_cp_element_group_909: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_909"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(907) & zeropad3D_CP_2067_elements(908);
      gj_zeropad3D_cp_element_group_909 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(909), clk => clk, reset => reset); --
    end block;
    -- CP-element group 910:  transition  input  bypass 
    -- CP-element group 910: predecessors 
    -- CP-element group 910: 	3 
    -- CP-element group 910: successors 
    -- CP-element group 910: 	912 
    -- CP-element group 910:  members (2) 
      -- CP-element group 910: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Sample/ra
      -- CP-element group 910: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Sample/$exit
      -- 
    ra_11505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 910_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_0, ack => zeropad3D_CP_2067_elements(910)); -- 
    -- CP-element group 911:  transition  input  bypass 
    -- CP-element group 911: predecessors 
    -- CP-element group 911: 	3 
    -- CP-element group 911: successors 
    -- CP-element group 911: 	912 
    -- CP-element group 911:  members (2) 
      -- CP-element group 911: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Update/ca
      -- CP-element group 911: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Update/$exit
      -- 
    ca_11510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 911_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_1, ack => zeropad3D_CP_2067_elements(911)); -- 
    -- CP-element group 912:  join  transition  output  bypass 
    -- CP-element group 912: predecessors 
    -- CP-element group 912: 	910 
    -- CP-element group 912: 	911 
    -- CP-element group 912: successors 
    -- CP-element group 912: 	916 
    -- CP-element group 912:  members (5) 
      -- CP-element group 912: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/$exit
      -- CP-element group 912: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_req
      -- CP-element group 912: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/$exit
      -- CP-element group 912: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/$exit
      -- CP-element group 912: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1797/$exit
      -- 
    phi_stmt_1797_req_11511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1797_req_11511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(912), ack => phi_stmt_1797_req_1); -- 
    zeropad3D_cp_element_group_912: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_912"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(910) & zeropad3D_CP_2067_elements(911);
      gj_zeropad3D_cp_element_group_912 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(912), clk => clk, reset => reset); --
    end block;
    -- CP-element group 913:  transition  input  bypass 
    -- CP-element group 913: predecessors 
    -- CP-element group 913: 	3 
    -- CP-element group 913: successors 
    -- CP-element group 913: 	915 
    -- CP-element group 913:  members (2) 
      -- CP-element group 913: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Sample/ra
      -- CP-element group 913: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Sample/$exit
      -- 
    ra_11528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 913_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1793_inst_ack_0, ack => zeropad3D_CP_2067_elements(913)); -- 
    -- CP-element group 914:  transition  input  bypass 
    -- CP-element group 914: predecessors 
    -- CP-element group 914: 	3 
    -- CP-element group 914: successors 
    -- CP-element group 914: 	915 
    -- CP-element group 914:  members (2) 
      -- CP-element group 914: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Update/$exit
      -- CP-element group 914: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Update/ca
      -- 
    ca_11533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 914_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1793_inst_ack_1, ack => zeropad3D_CP_2067_elements(914)); -- 
    -- CP-element group 915:  join  transition  output  bypass 
    -- CP-element group 915: predecessors 
    -- CP-element group 915: 	913 
    -- CP-element group 915: 	914 
    -- CP-element group 915: successors 
    -- CP-element group 915: 	916 
    -- CP-element group 915:  members (5) 
      -- CP-element group 915: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_req
      -- CP-element group 915: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/$exit
      -- CP-element group 915: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/$exit
      -- CP-element group 915: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/$exit
      -- CP-element group 915: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/phi_stmt_1790/$exit
      -- 
    phi_stmt_1790_req_11534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1790_req_11534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(915), ack => phi_stmt_1790_req_0); -- 
    zeropad3D_cp_element_group_915: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_915"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(913) & zeropad3D_CP_2067_elements(914);
      gj_zeropad3D_cp_element_group_915 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(915), clk => clk, reset => reset); --
    end block;
    -- CP-element group 916:  join  transition  bypass 
    -- CP-element group 916: predecessors 
    -- CP-element group 916: 	909 
    -- CP-element group 916: 	912 
    -- CP-element group 916: 	915 
    -- CP-element group 916: successors 
    -- CP-element group 916: 	923 
    -- CP-element group 916:  members (1) 
      -- CP-element group 916: 	 branch_block_stmt_655/ifx_xend607_whilex_xbody450_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_916: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_916"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(909) & zeropad3D_CP_2067_elements(912) & zeropad3D_CP_2067_elements(915);
      gj_zeropad3D_cp_element_group_916 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(916), clk => clk, reset => reset); --
    end block;
    -- CP-element group 917:  transition  output  delay-element  bypass 
    -- CP-element group 917: predecessors 
    -- CP-element group 917: 	227 
    -- CP-element group 917: successors 
    -- CP-element group 917: 	922 
    -- CP-element group 917:  members (4) 
      -- CP-element group 917: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_req
      -- CP-element group 917: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1807_konst_delay_trans
      -- CP-element group 917: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$exit
      -- CP-element group 917: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1803/$exit
      -- 
    phi_stmt_1803_req_11545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1803_req_11545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(917), ack => phi_stmt_1803_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(917) is a control-delay.
    cp_element_917_delay: control_delay_element  generic map(name => " 917_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(227), ack => zeropad3D_CP_2067_elements(917), clk => clk, reset =>reset);
    -- CP-element group 918:  transition  input  bypass 
    -- CP-element group 918: predecessors 
    -- CP-element group 918: 	227 
    -- CP-element group 918: successors 
    -- CP-element group 918: 	920 
    -- CP-element group 918:  members (2) 
      -- CP-element group 918: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Sample/ra
      -- CP-element group 918: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Sample/$exit
      -- 
    ra_11562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 918_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1800_inst_ack_0, ack => zeropad3D_CP_2067_elements(918)); -- 
    -- CP-element group 919:  transition  input  bypass 
    -- CP-element group 919: predecessors 
    -- CP-element group 919: 	227 
    -- CP-element group 919: successors 
    -- CP-element group 919: 	920 
    -- CP-element group 919:  members (2) 
      -- CP-element group 919: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Update/ca
      -- CP-element group 919: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Update/$exit
      -- 
    ca_11567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 919_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1800_inst_ack_1, ack => zeropad3D_CP_2067_elements(919)); -- 
    -- CP-element group 920:  join  transition  output  bypass 
    -- CP-element group 920: predecessors 
    -- CP-element group 920: 	918 
    -- CP-element group 920: 	919 
    -- CP-element group 920: successors 
    -- CP-element group 920: 	922 
    -- CP-element group 920:  members (5) 
      -- CP-element group 920: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/$exit
      -- CP-element group 920: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_req
      -- CP-element group 920: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/$exit
      -- CP-element group 920: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/$exit
      -- CP-element group 920: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/$exit
      -- 
    phi_stmt_1797_req_11568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1797_req_11568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(920), ack => phi_stmt_1797_req_0); -- 
    zeropad3D_cp_element_group_920: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_920"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(918) & zeropad3D_CP_2067_elements(919);
      gj_zeropad3D_cp_element_group_920 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(920), clk => clk, reset => reset); --
    end block;
    -- CP-element group 921:  transition  output  delay-element  bypass 
    -- CP-element group 921: predecessors 
    -- CP-element group 921: 	227 
    -- CP-element group 921: successors 
    -- CP-element group 921: 	922 
    -- CP-element group 921:  members (4) 
      -- CP-element group 921: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1790/$exit
      -- CP-element group 921: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/$exit
      -- CP-element group 921: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1796_konst_delay_trans
      -- CP-element group 921: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/phi_stmt_1790/phi_stmt_1790_req
      -- 
    phi_stmt_1790_req_11576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1790_req_11576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(921), ack => phi_stmt_1790_req_1); -- 
    -- Element group zeropad3D_CP_2067_elements(921) is a control-delay.
    cp_element_921_delay: control_delay_element  generic map(name => " 921_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(227), ack => zeropad3D_CP_2067_elements(921), clk => clk, reset =>reset);
    -- CP-element group 922:  join  transition  bypass 
    -- CP-element group 922: predecessors 
    -- CP-element group 922: 	917 
    -- CP-element group 922: 	920 
    -- CP-element group 922: 	921 
    -- CP-element group 922: successors 
    -- CP-element group 922: 	923 
    -- CP-element group 922:  members (1) 
      -- CP-element group 922: 	 branch_block_stmt_655/whilex_xend390_whilex_xbody450_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_922: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_922"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(917) & zeropad3D_CP_2067_elements(920) & zeropad3D_CP_2067_elements(921);
      gj_zeropad3D_cp_element_group_922 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(922), clk => clk, reset => reset); --
    end block;
    -- CP-element group 923:  merge  fork  transition  place  bypass 
    -- CP-element group 923: predecessors 
    -- CP-element group 923: 	916 
    -- CP-element group 923: 	922 
    -- CP-element group 923: successors 
    -- CP-element group 923: 	924 
    -- CP-element group 923: 	925 
    -- CP-element group 923: 	926 
    -- CP-element group 923:  members (2) 
      -- CP-element group 923: 	 branch_block_stmt_655/merge_stmt_1789_PhiReqMerge
      -- CP-element group 923: 	 branch_block_stmt_655/merge_stmt_1789_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(923) <= OrReduce(zeropad3D_CP_2067_elements(916) & zeropad3D_CP_2067_elements(922));
    -- CP-element group 924:  transition  input  bypass 
    -- CP-element group 924: predecessors 
    -- CP-element group 924: 	923 
    -- CP-element group 924: successors 
    -- CP-element group 924: 	927 
    -- CP-element group 924:  members (1) 
      -- CP-element group 924: 	 branch_block_stmt_655/merge_stmt_1789_PhiAck/phi_stmt_1790_ack
      -- 
    phi_stmt_1790_ack_11581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 924_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1790_ack_0, ack => zeropad3D_CP_2067_elements(924)); -- 
    -- CP-element group 925:  transition  input  bypass 
    -- CP-element group 925: predecessors 
    -- CP-element group 925: 	923 
    -- CP-element group 925: successors 
    -- CP-element group 925: 	927 
    -- CP-element group 925:  members (1) 
      -- CP-element group 925: 	 branch_block_stmt_655/merge_stmt_1789_PhiAck/phi_stmt_1797_ack
      -- 
    phi_stmt_1797_ack_11582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 925_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1797_ack_0, ack => zeropad3D_CP_2067_elements(925)); -- 
    -- CP-element group 926:  transition  input  bypass 
    -- CP-element group 926: predecessors 
    -- CP-element group 926: 	923 
    -- CP-element group 926: successors 
    -- CP-element group 926: 	927 
    -- CP-element group 926:  members (1) 
      -- CP-element group 926: 	 branch_block_stmt_655/merge_stmt_1789_PhiAck/phi_stmt_1803_ack
      -- 
    phi_stmt_1803_ack_11583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 926_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1803_ack_0, ack => zeropad3D_CP_2067_elements(926)); -- 
    -- CP-element group 927:  join  fork  transition  place  output  bypass 
    -- CP-element group 927: predecessors 
    -- CP-element group 927: 	924 
    -- CP-element group 927: 	925 
    -- CP-element group 927: 	926 
    -- CP-element group 927: successors 
    -- CP-element group 927: 	228 
    -- CP-element group 927: 	229 
    -- CP-element group 927:  members (10) 
      -- CP-element group 927: 	 branch_block_stmt_655/merge_stmt_1789__exit__
      -- CP-element group 927: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822__entry__
      -- CP-element group 927: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_Update/cr
      -- CP-element group 927: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_Update/$entry
      -- CP-element group 927: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_Sample/rr
      -- CP-element group 927: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_Sample/$entry
      -- CP-element group 927: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_update_start_
      -- CP-element group 927: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/type_cast_1814_sample_start_
      -- CP-element group 927: 	 branch_block_stmt_655/assign_stmt_1815_to_assign_stmt_1822/$entry
      -- CP-element group 927: 	 branch_block_stmt_655/merge_stmt_1789_PhiAck/$exit
      -- 
    cr_4805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(927), ack => type_cast_1814_inst_req_1); -- 
    rr_4800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(927), ack => type_cast_1814_inst_req_0); -- 
    zeropad3D_cp_element_group_927: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_927"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(924) & zeropad3D_CP_2067_elements(925) & zeropad3D_CP_2067_elements(926);
      gj_zeropad3D_cp_element_group_927 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(927), clk => clk, reset => reset); --
    end block;
    -- CP-element group 928:  merge  fork  transition  place  output  bypass 
    -- CP-element group 928: predecessors 
    -- CP-element group 928: 	230 
    -- CP-element group 928: 	237 
    -- CP-element group 928: 	240 
    -- CP-element group 928: 	247 
    -- CP-element group 928: successors 
    -- CP-element group 928: 	248 
    -- CP-element group 928: 	249 
    -- CP-element group 928: 	250 
    -- CP-element group 928: 	251 
    -- CP-element group 928: 	254 
    -- CP-element group 928: 	256 
    -- CP-element group 928: 	258 
    -- CP-element group 928: 	260 
    -- CP-element group 928:  members (33) 
      -- CP-element group 928: 	 branch_block_stmt_655/merge_stmt_1912__exit__
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968__entry__
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_sample_start_
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_update_start_
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_Sample/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_Sample/rr
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_Update/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1916_Update/cr
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_sample_start_
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_update_start_
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_Sample/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_Sample/rr
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_Update/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1921_Update/cr
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_update_start_
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_Update/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/type_cast_1955_Update/cr
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_update_start_
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_update_start
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_Update/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/array_obj_ref_1961_final_index_sum_regn_Update/req
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_complete/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/addr_of_1962_complete/req
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_update_start_
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Update/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Update/word_access_complete/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Update/word_access_complete/word_0/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/assign_stmt_1917_to_assign_stmt_1968/ptr_deref_1965_Update/word_access_complete/word_0/cr
      -- CP-element group 928: 	 branch_block_stmt_655/merge_stmt_1912_PhiReqMerge
      -- CP-element group 928: 	 branch_block_stmt_655/merge_stmt_1912_PhiAck/$entry
      -- CP-element group 928: 	 branch_block_stmt_655/merge_stmt_1912_PhiAck/$exit
      -- CP-element group 928: 	 branch_block_stmt_655/merge_stmt_1912_PhiAck/dummy
      -- 
    rr_5010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(928), ack => type_cast_1916_inst_req_0); -- 
    cr_5015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(928), ack => type_cast_1916_inst_req_1); -- 
    rr_5024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(928), ack => type_cast_1921_inst_req_0); -- 
    cr_5029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(928), ack => type_cast_1921_inst_req_1); -- 
    cr_5043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(928), ack => type_cast_1955_inst_req_1); -- 
    req_5074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(928), ack => array_obj_ref_1961_index_offset_req_1); -- 
    req_5089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(928), ack => addr_of_1962_final_reg_req_1); -- 
    cr_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(928), ack => ptr_deref_1965_store_0_req_1); -- 
    zeropad3D_CP_2067_elements(928) <= OrReduce(zeropad3D_CP_2067_elements(230) & zeropad3D_CP_2067_elements(237) & zeropad3D_CP_2067_elements(240) & zeropad3D_CP_2067_elements(247));
    -- CP-element group 929:  merge  fork  transition  place  output  bypass 
    -- CP-element group 929: predecessors 
    -- CP-element group 929: 	261 
    -- CP-element group 929: 	281 
    -- CP-element group 929: successors 
    -- CP-element group 929: 	282 
    -- CP-element group 929: 	283 
    -- CP-element group 929:  members (13) 
      -- CP-element group 929: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095__entry__
      -- CP-element group 929: 	 branch_block_stmt_655/merge_stmt_2077__exit__
      -- CP-element group 929: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/$entry
      -- CP-element group 929: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_sample_start_
      -- CP-element group 929: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_update_start_
      -- CP-element group 929: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_Sample/$entry
      -- CP-element group 929: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_Sample/rr
      -- CP-element group 929: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_Update/$entry
      -- CP-element group 929: 	 branch_block_stmt_655/assign_stmt_2082_to_assign_stmt_2095/type_cast_2081_Update/cr
      -- CP-element group 929: 	 branch_block_stmt_655/merge_stmt_2077_PhiReqMerge
      -- CP-element group 929: 	 branch_block_stmt_655/merge_stmt_2077_PhiAck/$entry
      -- CP-element group 929: 	 branch_block_stmt_655/merge_stmt_2077_PhiAck/$exit
      -- CP-element group 929: 	 branch_block_stmt_655/merge_stmt_2077_PhiAck/dummy
      -- 
    rr_5388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(929), ack => type_cast_2081_inst_req_0); -- 
    cr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(929), ack => type_cast_2081_inst_req_1); -- 
    zeropad3D_CP_2067_elements(929) <= OrReduce(zeropad3D_CP_2067_elements(261) & zeropad3D_CP_2067_elements(281));
    -- CP-element group 930:  transition  output  delay-element  bypass 
    -- CP-element group 930: predecessors 
    -- CP-element group 930: 	303 
    -- CP-element group 930: successors 
    -- CP-element group 930: 	937 
    -- CP-element group 930:  members (4) 
      -- CP-element group 930: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2196/$exit
      -- CP-element group 930: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/$exit
      -- CP-element group 930: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2202_konst_delay_trans
      -- CP-element group 930: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_req
      -- 
    phi_stmt_2196_req_11694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2196_req_11694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(930), ack => phi_stmt_2196_req_1); -- 
    -- Element group zeropad3D_CP_2067_elements(930) is a control-delay.
    cp_element_930_delay: control_delay_element  generic map(name => " 930_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(303), ack => zeropad3D_CP_2067_elements(930), clk => clk, reset =>reset);
    -- CP-element group 931:  transition  input  bypass 
    -- CP-element group 931: predecessors 
    -- CP-element group 931: 	303 
    -- CP-element group 931: successors 
    -- CP-element group 931: 	933 
    -- CP-element group 931:  members (2) 
      -- CP-element group 931: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/Sample/$exit
      -- CP-element group 931: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/Sample/ra
      -- 
    ra_11711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 931_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2206_inst_ack_0, ack => zeropad3D_CP_2067_elements(931)); -- 
    -- CP-element group 932:  transition  input  bypass 
    -- CP-element group 932: predecessors 
    -- CP-element group 932: 	303 
    -- CP-element group 932: successors 
    -- CP-element group 932: 	933 
    -- CP-element group 932:  members (2) 
      -- CP-element group 932: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/Update/$exit
      -- CP-element group 932: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/Update/ca
      -- 
    ca_11716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 932_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2206_inst_ack_1, ack => zeropad3D_CP_2067_elements(932)); -- 
    -- CP-element group 933:  join  transition  output  bypass 
    -- CP-element group 933: predecessors 
    -- CP-element group 933: 	931 
    -- CP-element group 933: 	932 
    -- CP-element group 933: successors 
    -- CP-element group 933: 	937 
    -- CP-element group 933:  members (5) 
      -- CP-element group 933: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/$exit
      -- CP-element group 933: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/$exit
      -- CP-element group 933: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/$exit
      -- CP-element group 933: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2206/SplitProtocol/$exit
      -- CP-element group 933: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_req
      -- 
    phi_stmt_2203_req_11717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2203_req_11717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(933), ack => phi_stmt_2203_req_0); -- 
    zeropad3D_cp_element_group_933: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_933"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(931) & zeropad3D_CP_2067_elements(932);
      gj_zeropad3D_cp_element_group_933 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(933), clk => clk, reset => reset); --
    end block;
    -- CP-element group 934:  transition  input  bypass 
    -- CP-element group 934: predecessors 
    -- CP-element group 934: 	303 
    -- CP-element group 934: successors 
    -- CP-element group 934: 	936 
    -- CP-element group 934:  members (2) 
      -- CP-element group 934: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/Sample/$exit
      -- CP-element group 934: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/Sample/ra
      -- 
    ra_11734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 934_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2212_inst_ack_0, ack => zeropad3D_CP_2067_elements(934)); -- 
    -- CP-element group 935:  transition  input  bypass 
    -- CP-element group 935: predecessors 
    -- CP-element group 935: 	303 
    -- CP-element group 935: successors 
    -- CP-element group 935: 	936 
    -- CP-element group 935:  members (2) 
      -- CP-element group 935: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/Update/$exit
      -- CP-element group 935: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/Update/ca
      -- 
    ca_11739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 935_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2212_inst_ack_1, ack => zeropad3D_CP_2067_elements(935)); -- 
    -- CP-element group 936:  join  transition  output  bypass 
    -- CP-element group 936: predecessors 
    -- CP-element group 936: 	934 
    -- CP-element group 936: 	935 
    -- CP-element group 936: successors 
    -- CP-element group 936: 	937 
    -- CP-element group 936:  members (5) 
      -- CP-element group 936: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/$exit
      -- CP-element group 936: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/$exit
      -- CP-element group 936: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/$exit
      -- CP-element group 936: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2212/SplitProtocol/$exit
      -- CP-element group 936: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_req
      -- 
    phi_stmt_2209_req_11740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2209_req_11740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(936), ack => phi_stmt_2209_req_0); -- 
    zeropad3D_cp_element_group_936: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_936"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(934) & zeropad3D_CP_2067_elements(935);
      gj_zeropad3D_cp_element_group_936 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(936), clk => clk, reset => reset); --
    end block;
    -- CP-element group 937:  join  transition  bypass 
    -- CP-element group 937: predecessors 
    -- CP-element group 937: 	930 
    -- CP-element group 937: 	933 
    -- CP-element group 937: 	936 
    -- CP-element group 937: successors 
    -- CP-element group 937: 	948 
    -- CP-element group 937:  members (1) 
      -- CP-element group 937: 	 branch_block_stmt_655/ifx_xelse570_ifx_xend607_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_937: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_937"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(930) & zeropad3D_CP_2067_elements(933) & zeropad3D_CP_2067_elements(936);
      gj_zeropad3D_cp_element_group_937 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(937), clk => clk, reset => reset); --
    end block;
    -- CP-element group 938:  transition  input  bypass 
    -- CP-element group 938: predecessors 
    -- CP-element group 938: 	284 
    -- CP-element group 938: successors 
    -- CP-element group 938: 	940 
    -- CP-element group 938:  members (2) 
      -- CP-element group 938: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/Sample/$exit
      -- CP-element group 938: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/Sample/ra
      -- 
    ra_11760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 938_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_0, ack => zeropad3D_CP_2067_elements(938)); -- 
    -- CP-element group 939:  transition  input  bypass 
    -- CP-element group 939: predecessors 
    -- CP-element group 939: 	284 
    -- CP-element group 939: successors 
    -- CP-element group 939: 	940 
    -- CP-element group 939:  members (2) 
      -- CP-element group 939: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/Update/$exit
      -- CP-element group 939: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/Update/ca
      -- 
    ca_11765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 939_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_1, ack => zeropad3D_CP_2067_elements(939)); -- 
    -- CP-element group 940:  join  transition  output  bypass 
    -- CP-element group 940: predecessors 
    -- CP-element group 940: 	938 
    -- CP-element group 940: 	939 
    -- CP-element group 940: successors 
    -- CP-element group 940: 	947 
    -- CP-element group 940:  members (5) 
      -- CP-element group 940: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/$exit
      -- CP-element group 940: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/$exit
      -- CP-element group 940: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/$exit
      -- CP-element group 940: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_sources/type_cast_2199/SplitProtocol/$exit
      -- CP-element group 940: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2196/phi_stmt_2196_req
      -- 
    phi_stmt_2196_req_11766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2196_req_11766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(940), ack => phi_stmt_2196_req_0); -- 
    zeropad3D_cp_element_group_940: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_940"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(938) & zeropad3D_CP_2067_elements(939);
      gj_zeropad3D_cp_element_group_940 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(940), clk => clk, reset => reset); --
    end block;
    -- CP-element group 941:  transition  input  bypass 
    -- CP-element group 941: predecessors 
    -- CP-element group 941: 	284 
    -- CP-element group 941: successors 
    -- CP-element group 941: 	943 
    -- CP-element group 941:  members (2) 
      -- CP-element group 941: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/Sample/$exit
      -- CP-element group 941: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/Sample/ra
      -- 
    ra_11783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 941_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2208_inst_ack_0, ack => zeropad3D_CP_2067_elements(941)); -- 
    -- CP-element group 942:  transition  input  bypass 
    -- CP-element group 942: predecessors 
    -- CP-element group 942: 	284 
    -- CP-element group 942: successors 
    -- CP-element group 942: 	943 
    -- CP-element group 942:  members (2) 
      -- CP-element group 942: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/Update/$exit
      -- CP-element group 942: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/Update/ca
      -- 
    ca_11788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 942_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2208_inst_ack_1, ack => zeropad3D_CP_2067_elements(942)); -- 
    -- CP-element group 943:  join  transition  output  bypass 
    -- CP-element group 943: predecessors 
    -- CP-element group 943: 	941 
    -- CP-element group 943: 	942 
    -- CP-element group 943: successors 
    -- CP-element group 943: 	947 
    -- CP-element group 943:  members (5) 
      -- CP-element group 943: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/$exit
      -- CP-element group 943: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/$exit
      -- CP-element group 943: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/$exit
      -- CP-element group 943: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_sources/type_cast_2208/SplitProtocol/$exit
      -- CP-element group 943: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2203/phi_stmt_2203_req
      -- 
    phi_stmt_2203_req_11789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2203_req_11789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(943), ack => phi_stmt_2203_req_1); -- 
    zeropad3D_cp_element_group_943: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_943"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(941) & zeropad3D_CP_2067_elements(942);
      gj_zeropad3D_cp_element_group_943 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(943), clk => clk, reset => reset); --
    end block;
    -- CP-element group 944:  transition  input  bypass 
    -- CP-element group 944: predecessors 
    -- CP-element group 944: 	284 
    -- CP-element group 944: successors 
    -- CP-element group 944: 	946 
    -- CP-element group 944:  members (2) 
      -- CP-element group 944: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/Sample/$exit
      -- CP-element group 944: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/Sample/ra
      -- 
    ra_11806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 944_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2214_inst_ack_0, ack => zeropad3D_CP_2067_elements(944)); -- 
    -- CP-element group 945:  transition  input  bypass 
    -- CP-element group 945: predecessors 
    -- CP-element group 945: 	284 
    -- CP-element group 945: successors 
    -- CP-element group 945: 	946 
    -- CP-element group 945:  members (2) 
      -- CP-element group 945: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/Update/$exit
      -- CP-element group 945: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/Update/ca
      -- 
    ca_11811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 945_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2214_inst_ack_1, ack => zeropad3D_CP_2067_elements(945)); -- 
    -- CP-element group 946:  join  transition  output  bypass 
    -- CP-element group 946: predecessors 
    -- CP-element group 946: 	944 
    -- CP-element group 946: 	945 
    -- CP-element group 946: successors 
    -- CP-element group 946: 	947 
    -- CP-element group 946:  members (5) 
      -- CP-element group 946: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/$exit
      -- CP-element group 946: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/$exit
      -- CP-element group 946: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/$exit
      -- CP-element group 946: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_sources/type_cast_2214/SplitProtocol/$exit
      -- CP-element group 946: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/phi_stmt_2209/phi_stmt_2209_req
      -- 
    phi_stmt_2209_req_11812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2209_req_11812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(946), ack => phi_stmt_2209_req_1); -- 
    zeropad3D_cp_element_group_946: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_946"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(944) & zeropad3D_CP_2067_elements(945);
      gj_zeropad3D_cp_element_group_946 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(946), clk => clk, reset => reset); --
    end block;
    -- CP-element group 947:  join  transition  bypass 
    -- CP-element group 947: predecessors 
    -- CP-element group 947: 	940 
    -- CP-element group 947: 	943 
    -- CP-element group 947: 	946 
    -- CP-element group 947: successors 
    -- CP-element group 947: 	948 
    -- CP-element group 947:  members (1) 
      -- CP-element group 947: 	 branch_block_stmt_655/ifx_xthen565_ifx_xend607_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_947: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_947"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(940) & zeropad3D_CP_2067_elements(943) & zeropad3D_CP_2067_elements(946);
      gj_zeropad3D_cp_element_group_947 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(947), clk => clk, reset => reset); --
    end block;
    -- CP-element group 948:  merge  fork  transition  place  bypass 
    -- CP-element group 948: predecessors 
    -- CP-element group 948: 	937 
    -- CP-element group 948: 	947 
    -- CP-element group 948: successors 
    -- CP-element group 948: 	949 
    -- CP-element group 948: 	950 
    -- CP-element group 948: 	951 
    -- CP-element group 948:  members (2) 
      -- CP-element group 948: 	 branch_block_stmt_655/merge_stmt_2195_PhiReqMerge
      -- CP-element group 948: 	 branch_block_stmt_655/merge_stmt_2195_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(948) <= OrReduce(zeropad3D_CP_2067_elements(937) & zeropad3D_CP_2067_elements(947));
    -- CP-element group 949:  transition  input  bypass 
    -- CP-element group 949: predecessors 
    -- CP-element group 949: 	948 
    -- CP-element group 949: successors 
    -- CP-element group 949: 	952 
    -- CP-element group 949:  members (1) 
      -- CP-element group 949: 	 branch_block_stmt_655/merge_stmt_2195_PhiAck/phi_stmt_2196_ack
      -- 
    phi_stmt_2196_ack_11817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 949_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2196_ack_0, ack => zeropad3D_CP_2067_elements(949)); -- 
    -- CP-element group 950:  transition  input  bypass 
    -- CP-element group 950: predecessors 
    -- CP-element group 950: 	948 
    -- CP-element group 950: successors 
    -- CP-element group 950: 	952 
    -- CP-element group 950:  members (1) 
      -- CP-element group 950: 	 branch_block_stmt_655/merge_stmt_2195_PhiAck/phi_stmt_2203_ack
      -- 
    phi_stmt_2203_ack_11818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 950_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2203_ack_0, ack => zeropad3D_CP_2067_elements(950)); -- 
    -- CP-element group 951:  transition  input  bypass 
    -- CP-element group 951: predecessors 
    -- CP-element group 951: 	948 
    -- CP-element group 951: successors 
    -- CP-element group 951: 	952 
    -- CP-element group 951:  members (1) 
      -- CP-element group 951: 	 branch_block_stmt_655/merge_stmt_2195_PhiAck/phi_stmt_2209_ack
      -- 
    phi_stmt_2209_ack_11819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 951_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2209_ack_0, ack => zeropad3D_CP_2067_elements(951)); -- 
    -- CP-element group 952:  join  transition  bypass 
    -- CP-element group 952: predecessors 
    -- CP-element group 952: 	949 
    -- CP-element group 952: 	950 
    -- CP-element group 952: 	951 
    -- CP-element group 952: successors 
    -- CP-element group 952: 	3 
    -- CP-element group 952:  members (1) 
      -- CP-element group 952: 	 branch_block_stmt_655/merge_stmt_2195_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_952: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_952"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(949) & zeropad3D_CP_2067_elements(950) & zeropad3D_CP_2067_elements(951);
      gj_zeropad3D_cp_element_group_952 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(952), clk => clk, reset => reset); --
    end block;
    -- CP-element group 953:  transition  input  bypass 
    -- CP-element group 953: predecessors 
    -- CP-element group 953: 	302 
    -- CP-element group 953: successors 
    -- CP-element group 953: 	955 
    -- CP-element group 953:  members (2) 
      -- CP-element group 953: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/Sample/$exit
      -- CP-element group 953: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/Sample/ra
      -- 
    ra_11839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 953_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2221_inst_ack_0, ack => zeropad3D_CP_2067_elements(953)); -- 
    -- CP-element group 954:  transition  input  bypass 
    -- CP-element group 954: predecessors 
    -- CP-element group 954: 	302 
    -- CP-element group 954: successors 
    -- CP-element group 954: 	955 
    -- CP-element group 954:  members (2) 
      -- CP-element group 954: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/Update/$exit
      -- CP-element group 954: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/Update/ca
      -- 
    ca_11844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 954_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2221_inst_ack_1, ack => zeropad3D_CP_2067_elements(954)); -- 
    -- CP-element group 955:  join  transition  output  bypass 
    -- CP-element group 955: predecessors 
    -- CP-element group 955: 	953 
    -- CP-element group 955: 	954 
    -- CP-element group 955: successors 
    -- CP-element group 955: 	962 
    -- CP-element group 955:  members (5) 
      -- CP-element group 955: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/$exit
      -- CP-element group 955: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/$exit
      -- CP-element group 955: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/$exit
      -- CP-element group 955: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_sources/type_cast_2221/SplitProtocol/$exit
      -- CP-element group 955: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2218/phi_stmt_2218_req
      -- 
    phi_stmt_2218_req_11845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2218_req_11845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(955), ack => phi_stmt_2218_req_0); -- 
    zeropad3D_cp_element_group_955: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_955"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(953) & zeropad3D_CP_2067_elements(954);
      gj_zeropad3D_cp_element_group_955 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(955), clk => clk, reset => reset); --
    end block;
    -- CP-element group 956:  transition  input  bypass 
    -- CP-element group 956: predecessors 
    -- CP-element group 956: 	302 
    -- CP-element group 956: successors 
    -- CP-element group 956: 	958 
    -- CP-element group 956:  members (2) 
      -- CP-element group 956: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/Sample/$exit
      -- CP-element group 956: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/Sample/ra
      -- 
    ra_11862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 956_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2225_inst_ack_0, ack => zeropad3D_CP_2067_elements(956)); -- 
    -- CP-element group 957:  transition  input  bypass 
    -- CP-element group 957: predecessors 
    -- CP-element group 957: 	302 
    -- CP-element group 957: successors 
    -- CP-element group 957: 	958 
    -- CP-element group 957:  members (2) 
      -- CP-element group 957: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/Update/$exit
      -- CP-element group 957: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/Update/ca
      -- 
    ca_11867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 957_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2225_inst_ack_1, ack => zeropad3D_CP_2067_elements(957)); -- 
    -- CP-element group 958:  join  transition  output  bypass 
    -- CP-element group 958: predecessors 
    -- CP-element group 958: 	956 
    -- CP-element group 958: 	957 
    -- CP-element group 958: successors 
    -- CP-element group 958: 	962 
    -- CP-element group 958:  members (5) 
      -- CP-element group 958: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/$exit
      -- CP-element group 958: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/$exit
      -- CP-element group 958: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/$exit
      -- CP-element group 958: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_sources/type_cast_2225/SplitProtocol/$exit
      -- CP-element group 958: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2222/phi_stmt_2222_req
      -- 
    phi_stmt_2222_req_11868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2222_req_11868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(958), ack => phi_stmt_2222_req_0); -- 
    zeropad3D_cp_element_group_958: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_958"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(956) & zeropad3D_CP_2067_elements(957);
      gj_zeropad3D_cp_element_group_958 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(958), clk => clk, reset => reset); --
    end block;
    -- CP-element group 959:  transition  input  bypass 
    -- CP-element group 959: predecessors 
    -- CP-element group 959: 	302 
    -- CP-element group 959: successors 
    -- CP-element group 959: 	961 
    -- CP-element group 959:  members (2) 
      -- CP-element group 959: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/Sample/$exit
      -- CP-element group 959: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/Sample/ra
      -- 
    ra_11885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 959_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2229_inst_ack_0, ack => zeropad3D_CP_2067_elements(959)); -- 
    -- CP-element group 960:  transition  input  bypass 
    -- CP-element group 960: predecessors 
    -- CP-element group 960: 	302 
    -- CP-element group 960: successors 
    -- CP-element group 960: 	961 
    -- CP-element group 960:  members (2) 
      -- CP-element group 960: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/Update/$exit
      -- CP-element group 960: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/Update/ca
      -- 
    ca_11890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 960_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2229_inst_ack_1, ack => zeropad3D_CP_2067_elements(960)); -- 
    -- CP-element group 961:  join  transition  output  bypass 
    -- CP-element group 961: predecessors 
    -- CP-element group 961: 	959 
    -- CP-element group 961: 	960 
    -- CP-element group 961: successors 
    -- CP-element group 961: 	962 
    -- CP-element group 961:  members (5) 
      -- CP-element group 961: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/$exit
      -- CP-element group 961: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/$exit
      -- CP-element group 961: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/$exit
      -- CP-element group 961: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_sources/type_cast_2229/SplitProtocol/$exit
      -- CP-element group 961: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/phi_stmt_2226/phi_stmt_2226_req
      -- 
    phi_stmt_2226_req_11891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2226_req_11891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(961), ack => phi_stmt_2226_req_0); -- 
    zeropad3D_cp_element_group_961: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_961"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(959) & zeropad3D_CP_2067_elements(960);
      gj_zeropad3D_cp_element_group_961 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(961), clk => clk, reset => reset); --
    end block;
    -- CP-element group 962:  join  fork  transition  place  bypass 
    -- CP-element group 962: predecessors 
    -- CP-element group 962: 	955 
    -- CP-element group 962: 	958 
    -- CP-element group 962: 	961 
    -- CP-element group 962: successors 
    -- CP-element group 962: 	963 
    -- CP-element group 962: 	964 
    -- CP-element group 962: 	965 
    -- CP-element group 962:  members (3) 
      -- CP-element group 962: 	 branch_block_stmt_655/ifx_xelse570_whilex_xend608_PhiReq/$exit
      -- CP-element group 962: 	 branch_block_stmt_655/merge_stmt_2217_PhiReqMerge
      -- CP-element group 962: 	 branch_block_stmt_655/merge_stmt_2217_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_962: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_962"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(955) & zeropad3D_CP_2067_elements(958) & zeropad3D_CP_2067_elements(961);
      gj_zeropad3D_cp_element_group_962 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(962), clk => clk, reset => reset); --
    end block;
    -- CP-element group 963:  transition  input  bypass 
    -- CP-element group 963: predecessors 
    -- CP-element group 963: 	962 
    -- CP-element group 963: successors 
    -- CP-element group 963: 	966 
    -- CP-element group 963:  members (1) 
      -- CP-element group 963: 	 branch_block_stmt_655/merge_stmt_2217_PhiAck/phi_stmt_2218_ack
      -- 
    phi_stmt_2218_ack_11896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 963_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2218_ack_0, ack => zeropad3D_CP_2067_elements(963)); -- 
    -- CP-element group 964:  transition  input  bypass 
    -- CP-element group 964: predecessors 
    -- CP-element group 964: 	962 
    -- CP-element group 964: successors 
    -- CP-element group 964: 	966 
    -- CP-element group 964:  members (1) 
      -- CP-element group 964: 	 branch_block_stmt_655/merge_stmt_2217_PhiAck/phi_stmt_2222_ack
      -- 
    phi_stmt_2222_ack_11897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 964_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2222_ack_0, ack => zeropad3D_CP_2067_elements(964)); -- 
    -- CP-element group 965:  transition  input  bypass 
    -- CP-element group 965: predecessors 
    -- CP-element group 965: 	962 
    -- CP-element group 965: successors 
    -- CP-element group 965: 	966 
    -- CP-element group 965:  members (1) 
      -- CP-element group 965: 	 branch_block_stmt_655/merge_stmt_2217_PhiAck/phi_stmt_2226_ack
      -- 
    phi_stmt_2226_ack_11898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 965_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2226_ack_0, ack => zeropad3D_CP_2067_elements(965)); -- 
    -- CP-element group 966:  join  fork  transition  place  output  bypass 
    -- CP-element group 966: predecessors 
    -- CP-element group 966: 	963 
    -- CP-element group 966: 	964 
    -- CP-element group 966: 	965 
    -- CP-element group 966: successors 
    -- CP-element group 966: 	304 
    -- CP-element group 966: 	305 
    -- CP-element group 966: 	306 
    -- CP-element group 966: 	307 
    -- CP-element group 966: 	308 
    -- CP-element group 966: 	309 
    -- CP-element group 966: 	310 
    -- CP-element group 966: 	311 
    -- CP-element group 966: 	312 
    -- CP-element group 966: 	313 
    -- CP-element group 966: 	314 
    -- CP-element group 966: 	315 
    -- CP-element group 966: 	317 
    -- CP-element group 966: 	319 
    -- CP-element group 966: 	321 
    -- CP-element group 966: 	323 
    -- CP-element group 966: 	325 
    -- CP-element group 966:  members (79) 
      -- CP-element group 966: 	 branch_block_stmt_655/merge_stmt_2217__exit__
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328__entry__
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_Update/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_Update/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2286_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_sample_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_Sample/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_Sample/rr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2233_Update/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_sample_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_Sample/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_Sample/rr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2243_Update/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_sample_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_word_address_calculated
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_root_address_calculated
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Sample/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Sample/word_access_start/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Sample/word_access_start/word_0/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Sample/word_access_start/word_0/rr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/word_access_complete/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/word_access_complete/word_0/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_pad_2252_Update/word_access_complete/word_0/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_sample_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_word_address_calculated
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_root_address_calculated
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Sample/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Sample/word_access_start/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Sample/word_access_start/word_0/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Sample/word_access_start/word_0/rr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/word_access_complete/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/word_access_complete/word_0/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_depth_high_2255_Update/word_access_complete/word_0/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_sample_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_word_address_calculated
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_root_address_calculated
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Sample/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Sample/word_access_start/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Sample/word_access_start/word_0/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Sample/word_access_start/word_0/rr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/word_access_complete/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/word_access_complete/word_0/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_depth_high_2258_Update/word_access_complete/word_0/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_sample_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_word_address_calculated
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_root_address_calculated
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Sample/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Sample/word_access_start/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Sample/word_access_start/word_0/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Sample/word_access_start/word_0/rr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/word_access_complete/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/word_access_complete/word_0/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/LOAD_out_col_high_2261_Update/word_access_complete/word_0/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2265_Update/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2269_Update/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_Update/$entry
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2273_Update/cr
      -- CP-element group 966: 	 branch_block_stmt_655/assign_stmt_2234_to_assign_stmt_2328/type_cast_2282_update_start_
      -- CP-element group 966: 	 branch_block_stmt_655/merge_stmt_2217_PhiAck/$exit
      -- 
    cr_5792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2282_inst_req_1); -- 
    cr_5806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2286_inst_req_1); -- 
    rr_5585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2233_inst_req_0); -- 
    cr_5590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2233_inst_req_1); -- 
    rr_5599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2243_inst_req_0); -- 
    cr_5604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2243_inst_req_1); -- 
    rr_5621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => LOAD_pad_2252_load_0_req_0); -- 
    cr_5632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => LOAD_pad_2252_load_0_req_1); -- 
    rr_5654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => LOAD_depth_high_2255_load_0_req_0); -- 
    cr_5665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => LOAD_depth_high_2255_load_0_req_1); -- 
    rr_5687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => LOAD_out_depth_high_2258_load_0_req_0); -- 
    cr_5698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => LOAD_out_depth_high_2258_load_0_req_1); -- 
    rr_5720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => LOAD_out_col_high_2261_load_0_req_0); -- 
    cr_5731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => LOAD_out_col_high_2261_load_0_req_1); -- 
    cr_5750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2265_inst_req_1); -- 
    cr_5764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2269_inst_req_1); -- 
    cr_5778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(966), ack => type_cast_2273_inst_req_1); -- 
    zeropad3D_cp_element_group_966: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_966"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(963) & zeropad3D_CP_2067_elements(964) & zeropad3D_CP_2067_elements(965);
      gj_zeropad3D_cp_element_group_966 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(966), clk => clk, reset => reset); --
    end block;
    -- CP-element group 967:  transition  input  bypass 
    -- CP-element group 967: predecessors 
    -- CP-element group 967: 	4 
    -- CP-element group 967: successors 
    -- CP-element group 967: 	969 
    -- CP-element group 967:  members (2) 
      -- CP-element group 967: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/Sample/$exit
      -- CP-element group 967: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/Sample/ra
      -- 
    ra_11918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 967_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2337_inst_ack_0, ack => zeropad3D_CP_2067_elements(967)); -- 
    -- CP-element group 968:  transition  input  bypass 
    -- CP-element group 968: predecessors 
    -- CP-element group 968: 	4 
    -- CP-element group 968: successors 
    -- CP-element group 968: 	969 
    -- CP-element group 968:  members (2) 
      -- CP-element group 968: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/Update/$exit
      -- CP-element group 968: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/Update/ca
      -- 
    ca_11923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 968_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2337_inst_ack_1, ack => zeropad3D_CP_2067_elements(968)); -- 
    -- CP-element group 969:  join  transition  output  bypass 
    -- CP-element group 969: predecessors 
    -- CP-element group 969: 	967 
    -- CP-element group 969: 	968 
    -- CP-element group 969: successors 
    -- CP-element group 969: 	976 
    -- CP-element group 969:  members (5) 
      -- CP-element group 969: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/$exit
      -- CP-element group 969: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/$exit
      -- CP-element group 969: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/$exit
      -- CP-element group 969: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2337/SplitProtocol/$exit
      -- CP-element group 969: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_req
      -- 
    phi_stmt_2331_req_11924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2331_req_11924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(969), ack => phi_stmt_2331_req_1); -- 
    zeropad3D_cp_element_group_969: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_969"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(967) & zeropad3D_CP_2067_elements(968);
      gj_zeropad3D_cp_element_group_969 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(969), clk => clk, reset => reset); --
    end block;
    -- CP-element group 970:  transition  input  bypass 
    -- CP-element group 970: predecessors 
    -- CP-element group 970: 	4 
    -- CP-element group 970: successors 
    -- CP-element group 970: 	972 
    -- CP-element group 970:  members (2) 
      -- CP-element group 970: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/Sample/$exit
      -- CP-element group 970: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/Sample/ra
      -- 
    ra_11941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 970_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2343_inst_ack_0, ack => zeropad3D_CP_2067_elements(970)); -- 
    -- CP-element group 971:  transition  input  bypass 
    -- CP-element group 971: predecessors 
    -- CP-element group 971: 	4 
    -- CP-element group 971: successors 
    -- CP-element group 971: 	972 
    -- CP-element group 971:  members (2) 
      -- CP-element group 971: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/Update/$exit
      -- CP-element group 971: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/Update/ca
      -- 
    ca_11946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 971_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2343_inst_ack_1, ack => zeropad3D_CP_2067_elements(971)); -- 
    -- CP-element group 972:  join  transition  output  bypass 
    -- CP-element group 972: predecessors 
    -- CP-element group 972: 	970 
    -- CP-element group 972: 	971 
    -- CP-element group 972: successors 
    -- CP-element group 972: 	976 
    -- CP-element group 972:  members (5) 
      -- CP-element group 972: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/$exit
      -- CP-element group 972: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/$exit
      -- CP-element group 972: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/$exit
      -- CP-element group 972: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2343/SplitProtocol/$exit
      -- CP-element group 972: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_req
      -- 
    phi_stmt_2338_req_11947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2338_req_11947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(972), ack => phi_stmt_2338_req_1); -- 
    zeropad3D_cp_element_group_972: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_972"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(970) & zeropad3D_CP_2067_elements(971);
      gj_zeropad3D_cp_element_group_972 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(972), clk => clk, reset => reset); --
    end block;
    -- CP-element group 973:  transition  input  bypass 
    -- CP-element group 973: predecessors 
    -- CP-element group 973: 	4 
    -- CP-element group 973: successors 
    -- CP-element group 973: 	975 
    -- CP-element group 973:  members (2) 
      -- CP-element group 973: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/Sample/$exit
      -- CP-element group 973: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/Sample/ra
      -- 
    ra_11964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 973_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2349_inst_ack_0, ack => zeropad3D_CP_2067_elements(973)); -- 
    -- CP-element group 974:  transition  input  bypass 
    -- CP-element group 974: predecessors 
    -- CP-element group 974: 	4 
    -- CP-element group 974: successors 
    -- CP-element group 974: 	975 
    -- CP-element group 974:  members (2) 
      -- CP-element group 974: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/Update/$exit
      -- CP-element group 974: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/Update/ca
      -- 
    ca_11969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 974_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2349_inst_ack_1, ack => zeropad3D_CP_2067_elements(974)); -- 
    -- CP-element group 975:  join  transition  output  bypass 
    -- CP-element group 975: predecessors 
    -- CP-element group 975: 	973 
    -- CP-element group 975: 	974 
    -- CP-element group 975: successors 
    -- CP-element group 975: 	976 
    -- CP-element group 975:  members (5) 
      -- CP-element group 975: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/$exit
      -- CP-element group 975: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/$exit
      -- CP-element group 975: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/$exit
      -- CP-element group 975: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2349/SplitProtocol/$exit
      -- CP-element group 975: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_req
      -- 
    phi_stmt_2344_req_11970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2344_req_11970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(975), ack => phi_stmt_2344_req_1); -- 
    zeropad3D_cp_element_group_975: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_975"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(973) & zeropad3D_CP_2067_elements(974);
      gj_zeropad3D_cp_element_group_975 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(975), clk => clk, reset => reset); --
    end block;
    -- CP-element group 976:  join  transition  bypass 
    -- CP-element group 976: predecessors 
    -- CP-element group 976: 	969 
    -- CP-element group 976: 	972 
    -- CP-element group 976: 	975 
    -- CP-element group 976: successors 
    -- CP-element group 976: 	985 
    -- CP-element group 976:  members (1) 
      -- CP-element group 976: 	 branch_block_stmt_655/ifx_xend827_whilex_xbody672_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_976: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_976"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(969) & zeropad3D_CP_2067_elements(972) & zeropad3D_CP_2067_elements(975);
      gj_zeropad3D_cp_element_group_976 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(976), clk => clk, reset => reset); --
    end block;
    -- CP-element group 977:  transition  output  delay-element  bypass 
    -- CP-element group 977: predecessors 
    -- CP-element group 977: 	326 
    -- CP-element group 977: successors 
    -- CP-element group 977: 	984 
    -- CP-element group 977:  members (4) 
      -- CP-element group 977: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2331/$exit
      -- CP-element group 977: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/$exit
      -- CP-element group 977: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_sources/type_cast_2335_konst_delay_trans
      -- CP-element group 977: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2331/phi_stmt_2331_req
      -- 
    phi_stmt_2331_req_11981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2331_req_11981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(977), ack => phi_stmt_2331_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(977) is a control-delay.
    cp_element_977_delay: control_delay_element  generic map(name => " 977_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(326), ack => zeropad3D_CP_2067_elements(977), clk => clk, reset =>reset);
    -- CP-element group 978:  transition  input  bypass 
    -- CP-element group 978: predecessors 
    -- CP-element group 978: 	326 
    -- CP-element group 978: successors 
    -- CP-element group 978: 	980 
    -- CP-element group 978:  members (2) 
      -- CP-element group 978: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/Sample/$exit
      -- CP-element group 978: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/Sample/ra
      -- 
    ra_11998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 978_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_0, ack => zeropad3D_CP_2067_elements(978)); -- 
    -- CP-element group 979:  transition  input  bypass 
    -- CP-element group 979: predecessors 
    -- CP-element group 979: 	326 
    -- CP-element group 979: successors 
    -- CP-element group 979: 	980 
    -- CP-element group 979:  members (2) 
      -- CP-element group 979: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/Update/$exit
      -- CP-element group 979: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/Update/ca
      -- 
    ca_12003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 979_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_1, ack => zeropad3D_CP_2067_elements(979)); -- 
    -- CP-element group 980:  join  transition  output  bypass 
    -- CP-element group 980: predecessors 
    -- CP-element group 980: 	978 
    -- CP-element group 980: 	979 
    -- CP-element group 980: successors 
    -- CP-element group 980: 	984 
    -- CP-element group 980:  members (5) 
      -- CP-element group 980: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/$exit
      -- CP-element group 980: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/$exit
      -- CP-element group 980: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/$exit
      -- CP-element group 980: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_sources/type_cast_2341/SplitProtocol/$exit
      -- CP-element group 980: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2338/phi_stmt_2338_req
      -- 
    phi_stmt_2338_req_12004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2338_req_12004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(980), ack => phi_stmt_2338_req_0); -- 
    zeropad3D_cp_element_group_980: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_980"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(978) & zeropad3D_CP_2067_elements(979);
      gj_zeropad3D_cp_element_group_980 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(980), clk => clk, reset => reset); --
    end block;
    -- CP-element group 981:  transition  input  bypass 
    -- CP-element group 981: predecessors 
    -- CP-element group 981: 	326 
    -- CP-element group 981: successors 
    -- CP-element group 981: 	983 
    -- CP-element group 981:  members (2) 
      -- CP-element group 981: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/Sample/$exit
      -- CP-element group 981: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/Sample/ra
      -- 
    ra_12021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 981_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_0, ack => zeropad3D_CP_2067_elements(981)); -- 
    -- CP-element group 982:  transition  input  bypass 
    -- CP-element group 982: predecessors 
    -- CP-element group 982: 	326 
    -- CP-element group 982: successors 
    -- CP-element group 982: 	983 
    -- CP-element group 982:  members (2) 
      -- CP-element group 982: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/Update/$exit
      -- CP-element group 982: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/Update/ca
      -- 
    ca_12026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 982_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_1, ack => zeropad3D_CP_2067_elements(982)); -- 
    -- CP-element group 983:  join  transition  output  bypass 
    -- CP-element group 983: predecessors 
    -- CP-element group 983: 	981 
    -- CP-element group 983: 	982 
    -- CP-element group 983: successors 
    -- CP-element group 983: 	984 
    -- CP-element group 983:  members (5) 
      -- CP-element group 983: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/$exit
      -- CP-element group 983: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/$exit
      -- CP-element group 983: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/$exit
      -- CP-element group 983: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_sources/type_cast_2347/SplitProtocol/$exit
      -- CP-element group 983: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/phi_stmt_2344/phi_stmt_2344_req
      -- 
    phi_stmt_2344_req_12027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2344_req_12027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(983), ack => phi_stmt_2344_req_0); -- 
    zeropad3D_cp_element_group_983: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_983"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(981) & zeropad3D_CP_2067_elements(982);
      gj_zeropad3D_cp_element_group_983 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(983), clk => clk, reset => reset); --
    end block;
    -- CP-element group 984:  join  transition  bypass 
    -- CP-element group 984: predecessors 
    -- CP-element group 984: 	977 
    -- CP-element group 984: 	980 
    -- CP-element group 984: 	983 
    -- CP-element group 984: successors 
    -- CP-element group 984: 	985 
    -- CP-element group 984:  members (1) 
      -- CP-element group 984: 	 branch_block_stmt_655/whilex_xend608_whilex_xbody672_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_984: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_984"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(977) & zeropad3D_CP_2067_elements(980) & zeropad3D_CP_2067_elements(983);
      gj_zeropad3D_cp_element_group_984 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(984), clk => clk, reset => reset); --
    end block;
    -- CP-element group 985:  merge  fork  transition  place  bypass 
    -- CP-element group 985: predecessors 
    -- CP-element group 985: 	976 
    -- CP-element group 985: 	984 
    -- CP-element group 985: successors 
    -- CP-element group 985: 	986 
    -- CP-element group 985: 	987 
    -- CP-element group 985: 	988 
    -- CP-element group 985:  members (2) 
      -- CP-element group 985: 	 branch_block_stmt_655/merge_stmt_2330_PhiReqMerge
      -- CP-element group 985: 	 branch_block_stmt_655/merge_stmt_2330_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(985) <= OrReduce(zeropad3D_CP_2067_elements(976) & zeropad3D_CP_2067_elements(984));
    -- CP-element group 986:  transition  input  bypass 
    -- CP-element group 986: predecessors 
    -- CP-element group 986: 	985 
    -- CP-element group 986: successors 
    -- CP-element group 986: 	989 
    -- CP-element group 986:  members (1) 
      -- CP-element group 986: 	 branch_block_stmt_655/merge_stmt_2330_PhiAck/phi_stmt_2331_ack
      -- 
    phi_stmt_2331_ack_12032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 986_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2331_ack_0, ack => zeropad3D_CP_2067_elements(986)); -- 
    -- CP-element group 987:  transition  input  bypass 
    -- CP-element group 987: predecessors 
    -- CP-element group 987: 	985 
    -- CP-element group 987: successors 
    -- CP-element group 987: 	989 
    -- CP-element group 987:  members (1) 
      -- CP-element group 987: 	 branch_block_stmt_655/merge_stmt_2330_PhiAck/phi_stmt_2338_ack
      -- 
    phi_stmt_2338_ack_12033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 987_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2338_ack_0, ack => zeropad3D_CP_2067_elements(987)); -- 
    -- CP-element group 988:  transition  input  bypass 
    -- CP-element group 988: predecessors 
    -- CP-element group 988: 	985 
    -- CP-element group 988: successors 
    -- CP-element group 988: 	989 
    -- CP-element group 988:  members (1) 
      -- CP-element group 988: 	 branch_block_stmt_655/merge_stmt_2330_PhiAck/phi_stmt_2344_ack
      -- 
    phi_stmt_2344_ack_12034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 988_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2344_ack_0, ack => zeropad3D_CP_2067_elements(988)); -- 
    -- CP-element group 989:  join  fork  transition  place  output  bypass 
    -- CP-element group 989: predecessors 
    -- CP-element group 989: 	986 
    -- CP-element group 989: 	987 
    -- CP-element group 989: 	988 
    -- CP-element group 989: successors 
    -- CP-element group 989: 	327 
    -- CP-element group 989: 	328 
    -- CP-element group 989:  members (10) 
      -- CP-element group 989: 	 branch_block_stmt_655/merge_stmt_2330__exit__
      -- CP-element group 989: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362__entry__
      -- CP-element group 989: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_update_start_
      -- CP-element group 989: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_Sample/$entry
      -- CP-element group 989: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_Update/cr
      -- CP-element group 989: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_sample_start_
      -- CP-element group 989: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/$entry
      -- CP-element group 989: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_Update/$entry
      -- CP-element group 989: 	 branch_block_stmt_655/assign_stmt_2355_to_assign_stmt_2362/type_cast_2354_Sample/rr
      -- CP-element group 989: 	 branch_block_stmt_655/merge_stmt_2330_PhiAck/$exit
      -- 
    cr_5823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(989), ack => type_cast_2354_inst_req_1); -- 
    rr_5818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(989), ack => type_cast_2354_inst_req_0); -- 
    zeropad3D_cp_element_group_989: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_989"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(986) & zeropad3D_CP_2067_elements(987) & zeropad3D_CP_2067_elements(988);
      gj_zeropad3D_cp_element_group_989 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(989), clk => clk, reset => reset); --
    end block;
    -- CP-element group 990:  merge  fork  transition  place  output  bypass 
    -- CP-element group 990: predecessors 
    -- CP-element group 990: 	329 
    -- CP-element group 990: 	336 
    -- CP-element group 990: 	339 
    -- CP-element group 990: 	346 
    -- CP-element group 990: successors 
    -- CP-element group 990: 	347 
    -- CP-element group 990: 	348 
    -- CP-element group 990: 	349 
    -- CP-element group 990: 	350 
    -- CP-element group 990: 	353 
    -- CP-element group 990: 	355 
    -- CP-element group 990: 	357 
    -- CP-element group 990: 	359 
    -- CP-element group 990:  members (33) 
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502__entry__
      -- CP-element group 990: 	 branch_block_stmt_655/merge_stmt_2446__exit__
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_sample_start_
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_update_start_
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_Sample/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_Sample/rr
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_Update/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2450_Update/cr
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_sample_start_
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_update_start_
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_Sample/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_Sample/rr
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_Update/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2455_Update/cr
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_update_start_
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_Update/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/type_cast_2489_Update/cr
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_update_start_
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_update_start
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_Update/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/array_obj_ref_2495_final_index_sum_regn_Update/req
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_complete/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/addr_of_2496_complete/req
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_update_start_
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Update/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Update/word_access_complete/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Update/word_access_complete/word_0/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/assign_stmt_2451_to_assign_stmt_2502/ptr_deref_2499_Update/word_access_complete/word_0/cr
      -- CP-element group 990: 	 branch_block_stmt_655/merge_stmt_2446_PhiReqMerge
      -- CP-element group 990: 	 branch_block_stmt_655/merge_stmt_2446_PhiAck/$entry
      -- CP-element group 990: 	 branch_block_stmt_655/merge_stmt_2446_PhiAck/$exit
      -- CP-element group 990: 	 branch_block_stmt_655/merge_stmt_2446_PhiAck/dummy
      -- 
    rr_6028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(990), ack => type_cast_2450_inst_req_0); -- 
    cr_6033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(990), ack => type_cast_2450_inst_req_1); -- 
    rr_6042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(990), ack => type_cast_2455_inst_req_0); -- 
    cr_6047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(990), ack => type_cast_2455_inst_req_1); -- 
    cr_6061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(990), ack => type_cast_2489_inst_req_1); -- 
    req_6092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(990), ack => array_obj_ref_2495_index_offset_req_1); -- 
    req_6107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(990), ack => addr_of_2496_final_reg_req_1); -- 
    cr_6157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(990), ack => ptr_deref_2499_store_0_req_1); -- 
    zeropad3D_CP_2067_elements(990) <= OrReduce(zeropad3D_CP_2067_elements(329) & zeropad3D_CP_2067_elements(336) & zeropad3D_CP_2067_elements(339) & zeropad3D_CP_2067_elements(346));
    -- CP-element group 991:  merge  fork  transition  place  output  bypass 
    -- CP-element group 991: predecessors 
    -- CP-element group 991: 	360 
    -- CP-element group 991: 	380 
    -- CP-element group 991: successors 
    -- CP-element group 991: 	381 
    -- CP-element group 991: 	382 
    -- CP-element group 991:  members (13) 
      -- CP-element group 991: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629__entry__
      -- CP-element group 991: 	 branch_block_stmt_655/merge_stmt_2611__exit__
      -- CP-element group 991: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/$entry
      -- CP-element group 991: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_sample_start_
      -- CP-element group 991: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_update_start_
      -- CP-element group 991: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_Sample/$entry
      -- CP-element group 991: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_Sample/rr
      -- CP-element group 991: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_Update/$entry
      -- CP-element group 991: 	 branch_block_stmt_655/assign_stmt_2616_to_assign_stmt_2629/type_cast_2615_Update/cr
      -- CP-element group 991: 	 branch_block_stmt_655/merge_stmt_2611_PhiReqMerge
      -- CP-element group 991: 	 branch_block_stmt_655/merge_stmt_2611_PhiAck/$entry
      -- CP-element group 991: 	 branch_block_stmt_655/merge_stmt_2611_PhiAck/$exit
      -- CP-element group 991: 	 branch_block_stmt_655/merge_stmt_2611_PhiAck/dummy
      -- 
    rr_6406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(991), ack => type_cast_2615_inst_req_0); -- 
    cr_6411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(991), ack => type_cast_2615_inst_req_1); -- 
    zeropad3D_CP_2067_elements(991) <= OrReduce(zeropad3D_CP_2067_elements(360) & zeropad3D_CP_2067_elements(380));
    -- CP-element group 992:  transition  output  delay-element  bypass 
    -- CP-element group 992: predecessors 
    -- CP-element group 992: 	402 
    -- CP-element group 992: successors 
    -- CP-element group 992: 	999 
    -- CP-element group 992:  members (4) 
      -- CP-element group 992: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2723/$exit
      -- CP-element group 992: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/$exit
      -- CP-element group 992: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2729_konst_delay_trans
      -- CP-element group 992: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_req
      -- 
    phi_stmt_2723_req_12145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2723_req_12145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(992), ack => phi_stmt_2723_req_1); -- 
    -- Element group zeropad3D_CP_2067_elements(992) is a control-delay.
    cp_element_992_delay: control_delay_element  generic map(name => " 992_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(402), ack => zeropad3D_CP_2067_elements(992), clk => clk, reset =>reset);
    -- CP-element group 993:  transition  input  bypass 
    -- CP-element group 993: predecessors 
    -- CP-element group 993: 	402 
    -- CP-element group 993: successors 
    -- CP-element group 993: 	995 
    -- CP-element group 993:  members (2) 
      -- CP-element group 993: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/Sample/$exit
      -- CP-element group 993: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/Sample/ra
      -- 
    ra_12162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 993_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2735_inst_ack_0, ack => zeropad3D_CP_2067_elements(993)); -- 
    -- CP-element group 994:  transition  input  bypass 
    -- CP-element group 994: predecessors 
    -- CP-element group 994: 	402 
    -- CP-element group 994: successors 
    -- CP-element group 994: 	995 
    -- CP-element group 994:  members (2) 
      -- CP-element group 994: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/Update/$exit
      -- CP-element group 994: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/Update/ca
      -- 
    ca_12167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 994_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2735_inst_ack_1, ack => zeropad3D_CP_2067_elements(994)); -- 
    -- CP-element group 995:  join  transition  output  bypass 
    -- CP-element group 995: predecessors 
    -- CP-element group 995: 	993 
    -- CP-element group 995: 	994 
    -- CP-element group 995: successors 
    -- CP-element group 995: 	999 
    -- CP-element group 995:  members (5) 
      -- CP-element group 995: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/$exit
      -- CP-element group 995: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/$exit
      -- CP-element group 995: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/$exit
      -- CP-element group 995: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2735/SplitProtocol/$exit
      -- CP-element group 995: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_req
      -- 
    phi_stmt_2730_req_12168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2730_req_12168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(995), ack => phi_stmt_2730_req_1); -- 
    zeropad3D_cp_element_group_995: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_995"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(993) & zeropad3D_CP_2067_elements(994);
      gj_zeropad3D_cp_element_group_995 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(995), clk => clk, reset => reset); --
    end block;
    -- CP-element group 996:  transition  input  bypass 
    -- CP-element group 996: predecessors 
    -- CP-element group 996: 	402 
    -- CP-element group 996: successors 
    -- CP-element group 996: 	998 
    -- CP-element group 996:  members (2) 
      -- CP-element group 996: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/Sample/$exit
      -- CP-element group 996: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/Sample/ra
      -- 
    ra_12185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 996_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2741_inst_ack_0, ack => zeropad3D_CP_2067_elements(996)); -- 
    -- CP-element group 997:  transition  input  bypass 
    -- CP-element group 997: predecessors 
    -- CP-element group 997: 	402 
    -- CP-element group 997: successors 
    -- CP-element group 997: 	998 
    -- CP-element group 997:  members (2) 
      -- CP-element group 997: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/Update/$exit
      -- CP-element group 997: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/Update/ca
      -- 
    ca_12190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 997_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2741_inst_ack_1, ack => zeropad3D_CP_2067_elements(997)); -- 
    -- CP-element group 998:  join  transition  output  bypass 
    -- CP-element group 998: predecessors 
    -- CP-element group 998: 	996 
    -- CP-element group 998: 	997 
    -- CP-element group 998: successors 
    -- CP-element group 998: 	999 
    -- CP-element group 998:  members (5) 
      -- CP-element group 998: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/$exit
      -- CP-element group 998: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/$exit
      -- CP-element group 998: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/$exit
      -- CP-element group 998: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2741/SplitProtocol/$exit
      -- CP-element group 998: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_req
      -- 
    phi_stmt_2736_req_12191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2736_req_12191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(998), ack => phi_stmt_2736_req_1); -- 
    zeropad3D_cp_element_group_998: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_998"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(996) & zeropad3D_CP_2067_elements(997);
      gj_zeropad3D_cp_element_group_998 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(998), clk => clk, reset => reset); --
    end block;
    -- CP-element group 999:  join  transition  bypass 
    -- CP-element group 999: predecessors 
    -- CP-element group 999: 	992 
    -- CP-element group 999: 	995 
    -- CP-element group 999: 	998 
    -- CP-element group 999: successors 
    -- CP-element group 999: 	1010 
    -- CP-element group 999:  members (1) 
      -- CP-element group 999: 	 branch_block_stmt_655/ifx_xelse791_ifx_xend827_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_999: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_999"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(992) & zeropad3D_CP_2067_elements(995) & zeropad3D_CP_2067_elements(998);
      gj_zeropad3D_cp_element_group_999 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(999), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1000:  transition  input  bypass 
    -- CP-element group 1000: predecessors 
    -- CP-element group 1000: 	383 
    -- CP-element group 1000: successors 
    -- CP-element group 1000: 	1002 
    -- CP-element group 1000:  members (2) 
      -- CP-element group 1000: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Sample/$exit
      -- CP-element group 1000: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Sample/ra
      -- 
    ra_12211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1000_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2726_inst_ack_0, ack => zeropad3D_CP_2067_elements(1000)); -- 
    -- CP-element group 1001:  transition  input  bypass 
    -- CP-element group 1001: predecessors 
    -- CP-element group 1001: 	383 
    -- CP-element group 1001: successors 
    -- CP-element group 1001: 	1002 
    -- CP-element group 1001:  members (2) 
      -- CP-element group 1001: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Update/$exit
      -- CP-element group 1001: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Update/ca
      -- 
    ca_12216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1001_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2726_inst_ack_1, ack => zeropad3D_CP_2067_elements(1001)); -- 
    -- CP-element group 1002:  join  transition  output  bypass 
    -- CP-element group 1002: predecessors 
    -- CP-element group 1002: 	1000 
    -- CP-element group 1002: 	1001 
    -- CP-element group 1002: successors 
    -- CP-element group 1002: 	1009 
    -- CP-element group 1002:  members (5) 
      -- CP-element group 1002: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/$exit
      -- CP-element group 1002: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/$exit
      -- CP-element group 1002: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/$exit
      -- CP-element group 1002: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/$exit
      -- CP-element group 1002: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2723/phi_stmt_2723_req
      -- 
    phi_stmt_2723_req_12217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2723_req_12217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1002), ack => phi_stmt_2723_req_0); -- 
    zeropad3D_cp_element_group_1002: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1002"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1000) & zeropad3D_CP_2067_elements(1001);
      gj_zeropad3D_cp_element_group_1002 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1002), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1003:  transition  input  bypass 
    -- CP-element group 1003: predecessors 
    -- CP-element group 1003: 	383 
    -- CP-element group 1003: successors 
    -- CP-element group 1003: 	1005 
    -- CP-element group 1003:  members (2) 
      -- CP-element group 1003: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/Sample/$exit
      -- CP-element group 1003: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/Sample/ra
      -- 
    ra_12234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1003_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2733_inst_ack_0, ack => zeropad3D_CP_2067_elements(1003)); -- 
    -- CP-element group 1004:  transition  input  bypass 
    -- CP-element group 1004: predecessors 
    -- CP-element group 1004: 	383 
    -- CP-element group 1004: successors 
    -- CP-element group 1004: 	1005 
    -- CP-element group 1004:  members (2) 
      -- CP-element group 1004: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/Update/$exit
      -- CP-element group 1004: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/Update/ca
      -- 
    ca_12239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1004_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2733_inst_ack_1, ack => zeropad3D_CP_2067_elements(1004)); -- 
    -- CP-element group 1005:  join  transition  output  bypass 
    -- CP-element group 1005: predecessors 
    -- CP-element group 1005: 	1003 
    -- CP-element group 1005: 	1004 
    -- CP-element group 1005: successors 
    -- CP-element group 1005: 	1009 
    -- CP-element group 1005:  members (5) 
      -- CP-element group 1005: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/$exit
      -- CP-element group 1005: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/$exit
      -- CP-element group 1005: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/$exit
      -- CP-element group 1005: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_sources/type_cast_2733/SplitProtocol/$exit
      -- CP-element group 1005: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2730/phi_stmt_2730_req
      -- 
    phi_stmt_2730_req_12240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2730_req_12240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1005), ack => phi_stmt_2730_req_0); -- 
    zeropad3D_cp_element_group_1005: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1005"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1003) & zeropad3D_CP_2067_elements(1004);
      gj_zeropad3D_cp_element_group_1005 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1005), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1006:  transition  input  bypass 
    -- CP-element group 1006: predecessors 
    -- CP-element group 1006: 	383 
    -- CP-element group 1006: successors 
    -- CP-element group 1006: 	1008 
    -- CP-element group 1006:  members (2) 
      -- CP-element group 1006: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/Sample/$exit
      -- CP-element group 1006: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/Sample/ra
      -- 
    ra_12257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1006_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2739_inst_ack_0, ack => zeropad3D_CP_2067_elements(1006)); -- 
    -- CP-element group 1007:  transition  input  bypass 
    -- CP-element group 1007: predecessors 
    -- CP-element group 1007: 	383 
    -- CP-element group 1007: successors 
    -- CP-element group 1007: 	1008 
    -- CP-element group 1007:  members (2) 
      -- CP-element group 1007: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/Update/$exit
      -- CP-element group 1007: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/Update/ca
      -- 
    ca_12262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1007_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2739_inst_ack_1, ack => zeropad3D_CP_2067_elements(1007)); -- 
    -- CP-element group 1008:  join  transition  output  bypass 
    -- CP-element group 1008: predecessors 
    -- CP-element group 1008: 	1006 
    -- CP-element group 1008: 	1007 
    -- CP-element group 1008: successors 
    -- CP-element group 1008: 	1009 
    -- CP-element group 1008:  members (5) 
      -- CP-element group 1008: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/$exit
      -- CP-element group 1008: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/$exit
      -- CP-element group 1008: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/$exit
      -- CP-element group 1008: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_sources/type_cast_2739/SplitProtocol/$exit
      -- CP-element group 1008: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/phi_stmt_2736/phi_stmt_2736_req
      -- 
    phi_stmt_2736_req_12263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2736_req_12263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1008), ack => phi_stmt_2736_req_0); -- 
    zeropad3D_cp_element_group_1008: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1008"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1006) & zeropad3D_CP_2067_elements(1007);
      gj_zeropad3D_cp_element_group_1008 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1008), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1009:  join  transition  bypass 
    -- CP-element group 1009: predecessors 
    -- CP-element group 1009: 	1002 
    -- CP-element group 1009: 	1005 
    -- CP-element group 1009: 	1008 
    -- CP-element group 1009: successors 
    -- CP-element group 1009: 	1010 
    -- CP-element group 1009:  members (1) 
      -- CP-element group 1009: 	 branch_block_stmt_655/ifx_xthen786_ifx_xend827_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1009: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1009"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1002) & zeropad3D_CP_2067_elements(1005) & zeropad3D_CP_2067_elements(1008);
      gj_zeropad3D_cp_element_group_1009 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1009), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1010:  merge  fork  transition  place  bypass 
    -- CP-element group 1010: predecessors 
    -- CP-element group 1010: 	999 
    -- CP-element group 1010: 	1009 
    -- CP-element group 1010: successors 
    -- CP-element group 1010: 	1011 
    -- CP-element group 1010: 	1012 
    -- CP-element group 1010: 	1013 
    -- CP-element group 1010:  members (2) 
      -- CP-element group 1010: 	 branch_block_stmt_655/merge_stmt_2722_PhiReqMerge
      -- CP-element group 1010: 	 branch_block_stmt_655/merge_stmt_2722_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1010) <= OrReduce(zeropad3D_CP_2067_elements(999) & zeropad3D_CP_2067_elements(1009));
    -- CP-element group 1011:  transition  input  bypass 
    -- CP-element group 1011: predecessors 
    -- CP-element group 1011: 	1010 
    -- CP-element group 1011: successors 
    -- CP-element group 1011: 	1014 
    -- CP-element group 1011:  members (1) 
      -- CP-element group 1011: 	 branch_block_stmt_655/merge_stmt_2722_PhiAck/phi_stmt_2723_ack
      -- 
    phi_stmt_2723_ack_12268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1011_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2723_ack_0, ack => zeropad3D_CP_2067_elements(1011)); -- 
    -- CP-element group 1012:  transition  input  bypass 
    -- CP-element group 1012: predecessors 
    -- CP-element group 1012: 	1010 
    -- CP-element group 1012: successors 
    -- CP-element group 1012: 	1014 
    -- CP-element group 1012:  members (1) 
      -- CP-element group 1012: 	 branch_block_stmt_655/merge_stmt_2722_PhiAck/phi_stmt_2730_ack
      -- 
    phi_stmt_2730_ack_12269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1012_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2730_ack_0, ack => zeropad3D_CP_2067_elements(1012)); -- 
    -- CP-element group 1013:  transition  input  bypass 
    -- CP-element group 1013: predecessors 
    -- CP-element group 1013: 	1010 
    -- CP-element group 1013: successors 
    -- CP-element group 1013: 	1014 
    -- CP-element group 1013:  members (1) 
      -- CP-element group 1013: 	 branch_block_stmt_655/merge_stmt_2722_PhiAck/phi_stmt_2736_ack
      -- 
    phi_stmt_2736_ack_12270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1013_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2736_ack_0, ack => zeropad3D_CP_2067_elements(1013)); -- 
    -- CP-element group 1014:  join  transition  bypass 
    -- CP-element group 1014: predecessors 
    -- CP-element group 1014: 	1011 
    -- CP-element group 1014: 	1012 
    -- CP-element group 1014: 	1013 
    -- CP-element group 1014: successors 
    -- CP-element group 1014: 	4 
    -- CP-element group 1014:  members (1) 
      -- CP-element group 1014: 	 branch_block_stmt_655/merge_stmt_2722_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1014: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1014"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1011) & zeropad3D_CP_2067_elements(1012) & zeropad3D_CP_2067_elements(1013);
      gj_zeropad3D_cp_element_group_1014 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1014), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1015:  transition  input  bypass 
    -- CP-element group 1015: predecessors 
    -- CP-element group 1015: 	401 
    -- CP-element group 1015: successors 
    -- CP-element group 1015: 	1017 
    -- CP-element group 1015:  members (2) 
      -- CP-element group 1015: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/Sample/$exit
      -- CP-element group 1015: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/Sample/ra
      -- 
    ra_12290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1015_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2748_inst_ack_0, ack => zeropad3D_CP_2067_elements(1015)); -- 
    -- CP-element group 1016:  transition  input  bypass 
    -- CP-element group 1016: predecessors 
    -- CP-element group 1016: 	401 
    -- CP-element group 1016: successors 
    -- CP-element group 1016: 	1017 
    -- CP-element group 1016:  members (2) 
      -- CP-element group 1016: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/Update/$exit
      -- CP-element group 1016: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/Update/ca
      -- 
    ca_12295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1016_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2748_inst_ack_1, ack => zeropad3D_CP_2067_elements(1016)); -- 
    -- CP-element group 1017:  join  transition  output  bypass 
    -- CP-element group 1017: predecessors 
    -- CP-element group 1017: 	1015 
    -- CP-element group 1017: 	1016 
    -- CP-element group 1017: successors 
    -- CP-element group 1017: 	1021 
    -- CP-element group 1017:  members (5) 
      -- CP-element group 1017: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/$exit
      -- CP-element group 1017: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/$exit
      -- CP-element group 1017: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/$exit
      -- CP-element group 1017: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_sources/type_cast_2748/SplitProtocol/$exit
      -- CP-element group 1017: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2745/phi_stmt_2745_req
      -- 
    phi_stmt_2745_req_12296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2745_req_12296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1017), ack => phi_stmt_2745_req_0); -- 
    zeropad3D_cp_element_group_1017: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1017"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1015) & zeropad3D_CP_2067_elements(1016);
      gj_zeropad3D_cp_element_group_1017 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1017), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1018:  transition  input  bypass 
    -- CP-element group 1018: predecessors 
    -- CP-element group 1018: 	401 
    -- CP-element group 1018: successors 
    -- CP-element group 1018: 	1020 
    -- CP-element group 1018:  members (2) 
      -- CP-element group 1018: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/Sample/$exit
      -- CP-element group 1018: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/Sample/ra
      -- 
    ra_12313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1018_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2752_inst_ack_0, ack => zeropad3D_CP_2067_elements(1018)); -- 
    -- CP-element group 1019:  transition  input  bypass 
    -- CP-element group 1019: predecessors 
    -- CP-element group 1019: 	401 
    -- CP-element group 1019: successors 
    -- CP-element group 1019: 	1020 
    -- CP-element group 1019:  members (2) 
      -- CP-element group 1019: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/Update/$exit
      -- CP-element group 1019: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/Update/ca
      -- 
    ca_12318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1019_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2752_inst_ack_1, ack => zeropad3D_CP_2067_elements(1019)); -- 
    -- CP-element group 1020:  join  transition  output  bypass 
    -- CP-element group 1020: predecessors 
    -- CP-element group 1020: 	1018 
    -- CP-element group 1020: 	1019 
    -- CP-element group 1020: successors 
    -- CP-element group 1020: 	1021 
    -- CP-element group 1020:  members (5) 
      -- CP-element group 1020: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/$exit
      -- CP-element group 1020: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/$exit
      -- CP-element group 1020: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/$exit
      -- CP-element group 1020: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_sources/type_cast_2752/SplitProtocol/$exit
      -- CP-element group 1020: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/phi_stmt_2749/phi_stmt_2749_req
      -- 
    phi_stmt_2749_req_12319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2749_req_12319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1020), ack => phi_stmt_2749_req_0); -- 
    zeropad3D_cp_element_group_1020: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1020"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1018) & zeropad3D_CP_2067_elements(1019);
      gj_zeropad3D_cp_element_group_1020 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1020), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1021:  join  fork  transition  place  bypass 
    -- CP-element group 1021: predecessors 
    -- CP-element group 1021: 	1017 
    -- CP-element group 1021: 	1020 
    -- CP-element group 1021: successors 
    -- CP-element group 1021: 	1022 
    -- CP-element group 1021: 	1023 
    -- CP-element group 1021:  members (3) 
      -- CP-element group 1021: 	 branch_block_stmt_655/ifx_xelse791_whilex_xend828_PhiReq/$exit
      -- CP-element group 1021: 	 branch_block_stmt_655/merge_stmt_2744_PhiReqMerge
      -- CP-element group 1021: 	 branch_block_stmt_655/merge_stmt_2744_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_1021: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1021"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1017) & zeropad3D_CP_2067_elements(1020);
      gj_zeropad3D_cp_element_group_1021 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1021), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1022:  transition  input  bypass 
    -- CP-element group 1022: predecessors 
    -- CP-element group 1022: 	1021 
    -- CP-element group 1022: successors 
    -- CP-element group 1022: 	1024 
    -- CP-element group 1022:  members (1) 
      -- CP-element group 1022: 	 branch_block_stmt_655/merge_stmt_2744_PhiAck/phi_stmt_2745_ack
      -- 
    phi_stmt_2745_ack_12324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1022_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2745_ack_0, ack => zeropad3D_CP_2067_elements(1022)); -- 
    -- CP-element group 1023:  transition  input  bypass 
    -- CP-element group 1023: predecessors 
    -- CP-element group 1023: 	1021 
    -- CP-element group 1023: successors 
    -- CP-element group 1023: 	1024 
    -- CP-element group 1023:  members (1) 
      -- CP-element group 1023: 	 branch_block_stmt_655/merge_stmt_2744_PhiAck/phi_stmt_2749_ack
      -- 
    phi_stmt_2749_ack_12325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1023_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2749_ack_0, ack => zeropad3D_CP_2067_elements(1023)); -- 
    -- CP-element group 1024:  join  fork  transition  place  output  bypass 
    -- CP-element group 1024: predecessors 
    -- CP-element group 1024: 	1022 
    -- CP-element group 1024: 	1023 
    -- CP-element group 1024: successors 
    -- CP-element group 1024: 	403 
    -- CP-element group 1024: 	404 
    -- CP-element group 1024: 	405 
    -- CP-element group 1024: 	406 
    -- CP-element group 1024: 	407 
    -- CP-element group 1024: 	408 
    -- CP-element group 1024: 	409 
    -- CP-element group 1024: 	410 
    -- CP-element group 1024: 	411 
    -- CP-element group 1024: 	412 
    -- CP-element group 1024: 	414 
    -- CP-element group 1024: 	416 
    -- CP-element group 1024: 	418 
    -- CP-element group 1024: 	420 
    -- CP-element group 1024: 	422 
    -- CP-element group 1024:  members (73) 
      -- CP-element group 1024: 	 branch_block_stmt_655/merge_stmt_2744__exit__
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841__entry__
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/word_access_complete/word_0/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_Update/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Sample/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/word_access_complete/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Sample/word_access_start/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/word_access_complete/word_0/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_sample_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Sample/word_access_start/word_0/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2795_Update/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_sample_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/word_access_complete/word_0/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/word_access_complete/word_0/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Sample/word_access_start/word_0/rr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_root_address_calculated
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_word_address_calculated
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_word_address_calculated
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_root_address_calculated
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Sample/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Sample/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2799_Update/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_root_address_calculated
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_word_address_calculated
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_sample_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/word_access_complete/word_0/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/word_access_complete/word_0/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2786_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/word_access_complete/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/word_access_complete/word_0/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/word_access_complete/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_Update/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Sample/word_access_start/word_0/rr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_depth_high_2771_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Sample/word_access_start/word_0/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_depth_high_2768_Sample/word_access_start/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Sample/word_access_start/word_0/rr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2782_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Sample/word_access_start/word_0/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_Update/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/word_access_complete/word_0/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/word_access_complete/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_out_col_high_2774_Sample/word_access_start/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2778_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_sample_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_Sample/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_Sample/rr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/type_cast_2756_Update/cr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_sample_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_word_address_calculated
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_root_address_calculated
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Sample/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Sample/word_access_start/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Sample/word_access_start/word_0/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Sample/word_access_start/word_0/rr
      -- CP-element group 1024: 	 branch_block_stmt_655/assign_stmt_2757_to_assign_stmt_2841/LOAD_pad_2765_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_655/merge_stmt_2744_PhiAck/$exit
      -- 
    cr_6782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => type_cast_2786_inst_req_1); -- 
    cr_6702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => LOAD_out_depth_high_2771_load_0_req_1); -- 
    cr_6796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => type_cast_2795_inst_req_1); -- 
    cr_6735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => LOAD_out_col_high_2774_load_0_req_1); -- 
    rr_6691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => LOAD_out_depth_high_2771_load_0_req_0); -- 
    cr_6810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => type_cast_2799_inst_req_1); -- 
    cr_6669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => LOAD_depth_high_2768_load_0_req_1); -- 
    cr_6636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => LOAD_pad_2765_load_0_req_1); -- 
    cr_6768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => type_cast_2782_inst_req_1); -- 
    rr_6658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => LOAD_depth_high_2768_load_0_req_0); -- 
    rr_6724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => LOAD_out_col_high_2774_load_0_req_0); -- 
    cr_6754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => type_cast_2778_inst_req_1); -- 
    rr_6603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => type_cast_2756_inst_req_0); -- 
    cr_6608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => type_cast_2756_inst_req_1); -- 
    rr_6625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1024), ack => LOAD_pad_2765_load_0_req_0); -- 
    zeropad3D_cp_element_group_1024: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1024"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1022) & zeropad3D_CP_2067_elements(1023);
      gj_zeropad3D_cp_element_group_1024 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1024), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1025:  transition  input  bypass 
    -- CP-element group 1025: predecessors 
    -- CP-element group 1025: 	5 
    -- CP-element group 1025: successors 
    -- CP-element group 1025: 	1027 
    -- CP-element group 1025:  members (2) 
      -- CP-element group 1025: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/Sample/$exit
      -- CP-element group 1025: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/Sample/ra
      -- 
    ra_12345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1025_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2850_inst_ack_0, ack => zeropad3D_CP_2067_elements(1025)); -- 
    -- CP-element group 1026:  transition  input  bypass 
    -- CP-element group 1026: predecessors 
    -- CP-element group 1026: 	5 
    -- CP-element group 1026: successors 
    -- CP-element group 1026: 	1027 
    -- CP-element group 1026:  members (2) 
      -- CP-element group 1026: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/Update/$exit
      -- CP-element group 1026: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/Update/ca
      -- 
    ca_12350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1026_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2850_inst_ack_1, ack => zeropad3D_CP_2067_elements(1026)); -- 
    -- CP-element group 1027:  join  transition  output  bypass 
    -- CP-element group 1027: predecessors 
    -- CP-element group 1027: 	1025 
    -- CP-element group 1027: 	1026 
    -- CP-element group 1027: successors 
    -- CP-element group 1027: 	1034 
    -- CP-element group 1027:  members (5) 
      -- CP-element group 1027: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/$exit
      -- CP-element group 1027: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/$exit
      -- CP-element group 1027: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/$exit
      -- CP-element group 1027: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2850/SplitProtocol/$exit
      -- CP-element group 1027: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_req
      -- 
    phi_stmt_2844_req_12351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2844_req_12351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1027), ack => phi_stmt_2844_req_1); -- 
    zeropad3D_cp_element_group_1027: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1027"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1025) & zeropad3D_CP_2067_elements(1026);
      gj_zeropad3D_cp_element_group_1027 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1027), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1028:  transition  input  bypass 
    -- CP-element group 1028: predecessors 
    -- CP-element group 1028: 	5 
    -- CP-element group 1028: successors 
    -- CP-element group 1028: 	1030 
    -- CP-element group 1028:  members (2) 
      -- CP-element group 1028: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/Sample/$exit
      -- CP-element group 1028: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/Sample/ra
      -- 
    ra_12368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1028_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2856_inst_ack_0, ack => zeropad3D_CP_2067_elements(1028)); -- 
    -- CP-element group 1029:  transition  input  bypass 
    -- CP-element group 1029: predecessors 
    -- CP-element group 1029: 	5 
    -- CP-element group 1029: successors 
    -- CP-element group 1029: 	1030 
    -- CP-element group 1029:  members (2) 
      -- CP-element group 1029: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/Update/$exit
      -- CP-element group 1029: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/Update/ca
      -- 
    ca_12373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1029_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2856_inst_ack_1, ack => zeropad3D_CP_2067_elements(1029)); -- 
    -- CP-element group 1030:  join  transition  output  bypass 
    -- CP-element group 1030: predecessors 
    -- CP-element group 1030: 	1028 
    -- CP-element group 1030: 	1029 
    -- CP-element group 1030: successors 
    -- CP-element group 1030: 	1034 
    -- CP-element group 1030:  members (5) 
      -- CP-element group 1030: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/$exit
      -- CP-element group 1030: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/$exit
      -- CP-element group 1030: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/$exit
      -- CP-element group 1030: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2856/SplitProtocol/$exit
      -- CP-element group 1030: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_req
      -- 
    phi_stmt_2851_req_12374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2851_req_12374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1030), ack => phi_stmt_2851_req_1); -- 
    zeropad3D_cp_element_group_1030: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1030"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1028) & zeropad3D_CP_2067_elements(1029);
      gj_zeropad3D_cp_element_group_1030 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1030), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1031:  transition  input  bypass 
    -- CP-element group 1031: predecessors 
    -- CP-element group 1031: 	5 
    -- CP-element group 1031: successors 
    -- CP-element group 1031: 	1033 
    -- CP-element group 1031:  members (2) 
      -- CP-element group 1031: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/Sample/$exit
      -- CP-element group 1031: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/Sample/ra
      -- 
    ra_12391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1031_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2863_inst_ack_0, ack => zeropad3D_CP_2067_elements(1031)); -- 
    -- CP-element group 1032:  transition  input  bypass 
    -- CP-element group 1032: predecessors 
    -- CP-element group 1032: 	5 
    -- CP-element group 1032: successors 
    -- CP-element group 1032: 	1033 
    -- CP-element group 1032:  members (2) 
      -- CP-element group 1032: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/Update/$exit
      -- CP-element group 1032: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/Update/ca
      -- 
    ca_12396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1032_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2863_inst_ack_1, ack => zeropad3D_CP_2067_elements(1032)); -- 
    -- CP-element group 1033:  join  transition  output  bypass 
    -- CP-element group 1033: predecessors 
    -- CP-element group 1033: 	1031 
    -- CP-element group 1033: 	1032 
    -- CP-element group 1033: successors 
    -- CP-element group 1033: 	1034 
    -- CP-element group 1033:  members (5) 
      -- CP-element group 1033: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/$exit
      -- CP-element group 1033: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/$exit
      -- CP-element group 1033: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/$exit
      -- CP-element group 1033: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2863/SplitProtocol/$exit
      -- CP-element group 1033: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_req
      -- 
    phi_stmt_2857_req_12397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2857_req_12397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1033), ack => phi_stmt_2857_req_1); -- 
    zeropad3D_cp_element_group_1033: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1033"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1031) & zeropad3D_CP_2067_elements(1032);
      gj_zeropad3D_cp_element_group_1033 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1033), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1034:  join  transition  bypass 
    -- CP-element group 1034: predecessors 
    -- CP-element group 1034: 	1027 
    -- CP-element group 1034: 	1030 
    -- CP-element group 1034: 	1033 
    -- CP-element group 1034: successors 
    -- CP-element group 1034: 	1041 
    -- CP-element group 1034:  members (1) 
      -- CP-element group 1034: 	 branch_block_stmt_655/ifx_xend1047_whilex_xbody888_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1034: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1034"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1027) & zeropad3D_CP_2067_elements(1030) & zeropad3D_CP_2067_elements(1033);
      gj_zeropad3D_cp_element_group_1034 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1034), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1035:  transition  output  delay-element  bypass 
    -- CP-element group 1035: predecessors 
    -- CP-element group 1035: 	423 
    -- CP-element group 1035: successors 
    -- CP-element group 1035: 	1040 
    -- CP-element group 1035:  members (4) 
      -- CP-element group 1035: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2844/$exit
      -- CP-element group 1035: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/$exit
      -- CP-element group 1035: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_sources/type_cast_2848_konst_delay_trans
      -- CP-element group 1035: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2844/phi_stmt_2844_req
      -- 
    phi_stmt_2844_req_12408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2844_req_12408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1035), ack => phi_stmt_2844_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(1035) is a control-delay.
    cp_element_1035_delay: control_delay_element  generic map(name => " 1035_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(423), ack => zeropad3D_CP_2067_elements(1035), clk => clk, reset =>reset);
    -- CP-element group 1036:  transition  input  bypass 
    -- CP-element group 1036: predecessors 
    -- CP-element group 1036: 	423 
    -- CP-element group 1036: successors 
    -- CP-element group 1036: 	1038 
    -- CP-element group 1036:  members (2) 
      -- CP-element group 1036: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/Sample/$exit
      -- CP-element group 1036: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/Sample/ra
      -- 
    ra_12425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1036_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2854_inst_ack_0, ack => zeropad3D_CP_2067_elements(1036)); -- 
    -- CP-element group 1037:  transition  input  bypass 
    -- CP-element group 1037: predecessors 
    -- CP-element group 1037: 	423 
    -- CP-element group 1037: successors 
    -- CP-element group 1037: 	1038 
    -- CP-element group 1037:  members (2) 
      -- CP-element group 1037: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/Update/$exit
      -- CP-element group 1037: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/Update/ca
      -- 
    ca_12430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1037_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2854_inst_ack_1, ack => zeropad3D_CP_2067_elements(1037)); -- 
    -- CP-element group 1038:  join  transition  output  bypass 
    -- CP-element group 1038: predecessors 
    -- CP-element group 1038: 	1036 
    -- CP-element group 1038: 	1037 
    -- CP-element group 1038: successors 
    -- CP-element group 1038: 	1040 
    -- CP-element group 1038:  members (5) 
      -- CP-element group 1038: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/$exit
      -- CP-element group 1038: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/$exit
      -- CP-element group 1038: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/$exit
      -- CP-element group 1038: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_sources/type_cast_2854/SplitProtocol/$exit
      -- CP-element group 1038: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2851/phi_stmt_2851_req
      -- 
    phi_stmt_2851_req_12431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2851_req_12431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1038), ack => phi_stmt_2851_req_0); -- 
    zeropad3D_cp_element_group_1038: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1038"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1036) & zeropad3D_CP_2067_elements(1037);
      gj_zeropad3D_cp_element_group_1038 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1038), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1039:  transition  output  delay-element  bypass 
    -- CP-element group 1039: predecessors 
    -- CP-element group 1039: 	423 
    -- CP-element group 1039: successors 
    -- CP-element group 1039: 	1040 
    -- CP-element group 1039:  members (4) 
      -- CP-element group 1039: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2857/$exit
      -- CP-element group 1039: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/$exit
      -- CP-element group 1039: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_sources/type_cast_2861_konst_delay_trans
      -- CP-element group 1039: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/phi_stmt_2857/phi_stmt_2857_req
      -- 
    phi_stmt_2857_req_12439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2857_req_12439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1039), ack => phi_stmt_2857_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(1039) is a control-delay.
    cp_element_1039_delay: control_delay_element  generic map(name => " 1039_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(423), ack => zeropad3D_CP_2067_elements(1039), clk => clk, reset =>reset);
    -- CP-element group 1040:  join  transition  bypass 
    -- CP-element group 1040: predecessors 
    -- CP-element group 1040: 	1035 
    -- CP-element group 1040: 	1038 
    -- CP-element group 1040: 	1039 
    -- CP-element group 1040: successors 
    -- CP-element group 1040: 	1041 
    -- CP-element group 1040:  members (1) 
      -- CP-element group 1040: 	 branch_block_stmt_655/whilex_xend828_whilex_xbody888_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1040: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1040"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1035) & zeropad3D_CP_2067_elements(1038) & zeropad3D_CP_2067_elements(1039);
      gj_zeropad3D_cp_element_group_1040 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1040), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1041:  merge  fork  transition  place  bypass 
    -- CP-element group 1041: predecessors 
    -- CP-element group 1041: 	1034 
    -- CP-element group 1041: 	1040 
    -- CP-element group 1041: successors 
    -- CP-element group 1041: 	1042 
    -- CP-element group 1041: 	1043 
    -- CP-element group 1041: 	1044 
    -- CP-element group 1041:  members (2) 
      -- CP-element group 1041: 	 branch_block_stmt_655/merge_stmt_2843_PhiReqMerge
      -- CP-element group 1041: 	 branch_block_stmt_655/merge_stmt_2843_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1041) <= OrReduce(zeropad3D_CP_2067_elements(1034) & zeropad3D_CP_2067_elements(1040));
    -- CP-element group 1042:  transition  input  bypass 
    -- CP-element group 1042: predecessors 
    -- CP-element group 1042: 	1041 
    -- CP-element group 1042: successors 
    -- CP-element group 1042: 	1045 
    -- CP-element group 1042:  members (1) 
      -- CP-element group 1042: 	 branch_block_stmt_655/merge_stmt_2843_PhiAck/phi_stmt_2844_ack
      -- 
    phi_stmt_2844_ack_12444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1042_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2844_ack_0, ack => zeropad3D_CP_2067_elements(1042)); -- 
    -- CP-element group 1043:  transition  input  bypass 
    -- CP-element group 1043: predecessors 
    -- CP-element group 1043: 	1041 
    -- CP-element group 1043: successors 
    -- CP-element group 1043: 	1045 
    -- CP-element group 1043:  members (1) 
      -- CP-element group 1043: 	 branch_block_stmt_655/merge_stmt_2843_PhiAck/phi_stmt_2851_ack
      -- 
    phi_stmt_2851_ack_12445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1043_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2851_ack_0, ack => zeropad3D_CP_2067_elements(1043)); -- 
    -- CP-element group 1044:  transition  input  bypass 
    -- CP-element group 1044: predecessors 
    -- CP-element group 1044: 	1041 
    -- CP-element group 1044: successors 
    -- CP-element group 1044: 	1045 
    -- CP-element group 1044:  members (1) 
      -- CP-element group 1044: 	 branch_block_stmt_655/merge_stmt_2843_PhiAck/phi_stmt_2857_ack
      -- 
    phi_stmt_2857_ack_12446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1044_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2857_ack_0, ack => zeropad3D_CP_2067_elements(1044)); -- 
    -- CP-element group 1045:  join  fork  transition  place  output  bypass 
    -- CP-element group 1045: predecessors 
    -- CP-element group 1045: 	1042 
    -- CP-element group 1045: 	1043 
    -- CP-element group 1045: 	1044 
    -- CP-element group 1045: successors 
    -- CP-element group 1045: 	424 
    -- CP-element group 1045: 	425 
    -- CP-element group 1045:  members (10) 
      -- CP-element group 1045: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876__entry__
      -- CP-element group 1045: 	 branch_block_stmt_655/merge_stmt_2843__exit__
      -- CP-element group 1045: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_Update/cr
      -- CP-element group 1045: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_Update/$entry
      -- CP-element group 1045: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_Sample/rr
      -- CP-element group 1045: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_Sample/$entry
      -- CP-element group 1045: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_update_start_
      -- CP-element group 1045: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/type_cast_2868_sample_start_
      -- CP-element group 1045: 	 branch_block_stmt_655/assign_stmt_2869_to_assign_stmt_2876/$entry
      -- CP-element group 1045: 	 branch_block_stmt_655/merge_stmt_2843_PhiAck/$exit
      -- 
    cr_6827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1045), ack => type_cast_2868_inst_req_1); -- 
    rr_6822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1045), ack => type_cast_2868_inst_req_0); -- 
    zeropad3D_cp_element_group_1045: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1045"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1042) & zeropad3D_CP_2067_elements(1043) & zeropad3D_CP_2067_elements(1044);
      gj_zeropad3D_cp_element_group_1045 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1045), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1046:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1046: predecessors 
    -- CP-element group 1046: 	426 
    -- CP-element group 1046: 	433 
    -- CP-element group 1046: 	436 
    -- CP-element group 1046: 	443 
    -- CP-element group 1046: successors 
    -- CP-element group 1046: 	444 
    -- CP-element group 1046: 	445 
    -- CP-element group 1046: 	446 
    -- CP-element group 1046: 	447 
    -- CP-element group 1046: 	450 
    -- CP-element group 1046: 	452 
    -- CP-element group 1046: 	454 
    -- CP-element group 1046: 	456 
    -- CP-element group 1046:  members (33) 
      -- CP-element group 1046: 	 branch_block_stmt_655/merge_stmt_2972__exit__
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028__entry__
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_update_start_
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_sample_start_
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_Update/cr
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_Update/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_sample_start_
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_Update/cr
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_Update/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_3015_update_start_
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_Sample/rr
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_Update/cr
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_Update/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_Sample/rr
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2981_Sample/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_Sample/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/type_cast_2976_update_start_
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_update_start_
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_update_start
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_Update/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/array_obj_ref_3021_final_index_sum_regn_Update/req
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_complete/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/addr_of_3022_complete/req
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_update_start_
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Update/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Update/word_access_complete/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Update/word_access_complete/word_0/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/assign_stmt_2977_to_assign_stmt_3028/ptr_deref_3025_Update/word_access_complete/word_0/cr
      -- CP-element group 1046: 	 branch_block_stmt_655/merge_stmt_2972_PhiReqMerge
      -- CP-element group 1046: 	 branch_block_stmt_655/merge_stmt_2972_PhiAck/$entry
      -- CP-element group 1046: 	 branch_block_stmt_655/merge_stmt_2972_PhiAck/$exit
      -- CP-element group 1046: 	 branch_block_stmt_655/merge_stmt_2972_PhiAck/dummy
      -- 
    cr_7065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1046), ack => type_cast_3015_inst_req_1); -- 
    cr_7037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1046), ack => type_cast_2976_inst_req_1); -- 
    rr_7032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1046), ack => type_cast_2976_inst_req_0); -- 
    cr_7051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1046), ack => type_cast_2981_inst_req_1); -- 
    rr_7046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1046), ack => type_cast_2981_inst_req_0); -- 
    req_7096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1046), ack => array_obj_ref_3021_index_offset_req_1); -- 
    req_7111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1046), ack => addr_of_3022_final_reg_req_1); -- 
    cr_7161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1046), ack => ptr_deref_3025_store_0_req_1); -- 
    zeropad3D_CP_2067_elements(1046) <= OrReduce(zeropad3D_CP_2067_elements(426) & zeropad3D_CP_2067_elements(433) & zeropad3D_CP_2067_elements(436) & zeropad3D_CP_2067_elements(443));
    -- CP-element group 1047:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1047: predecessors 
    -- CP-element group 1047: 	457 
    -- CP-element group 1047: 	477 
    -- CP-element group 1047: successors 
    -- CP-element group 1047: 	478 
    -- CP-element group 1047: 	479 
    -- CP-element group 1047:  members (13) 
      -- CP-element group 1047: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155__entry__
      -- CP-element group 1047: 	 branch_block_stmt_655/merge_stmt_3137__exit__
      -- CP-element group 1047: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/$entry
      -- CP-element group 1047: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_sample_start_
      -- CP-element group 1047: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_update_start_
      -- CP-element group 1047: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_Sample/$entry
      -- CP-element group 1047: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_Sample/rr
      -- CP-element group 1047: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_Update/$entry
      -- CP-element group 1047: 	 branch_block_stmt_655/assign_stmt_3142_to_assign_stmt_3155/type_cast_3141_Update/cr
      -- CP-element group 1047: 	 branch_block_stmt_655/merge_stmt_3137_PhiReqMerge
      -- CP-element group 1047: 	 branch_block_stmt_655/merge_stmt_3137_PhiAck/$entry
      -- CP-element group 1047: 	 branch_block_stmt_655/merge_stmt_3137_PhiAck/$exit
      -- CP-element group 1047: 	 branch_block_stmt_655/merge_stmt_3137_PhiAck/dummy
      -- 
    rr_7410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1047), ack => type_cast_3141_inst_req_0); -- 
    cr_7415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1047), ack => type_cast_3141_inst_req_1); -- 
    zeropad3D_CP_2067_elements(1047) <= OrReduce(zeropad3D_CP_2067_elements(457) & zeropad3D_CP_2067_elements(477));
    -- CP-element group 1048:  transition  input  bypass 
    -- CP-element group 1048: predecessors 
    -- CP-element group 1048: 	499 
    -- CP-element group 1048: successors 
    -- CP-element group 1048: 	1050 
    -- CP-element group 1048:  members (2) 
      -- CP-element group 1048: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/Sample/$exit
      -- CP-element group 1048: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/Sample/ra
      -- 
    ra_12566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1048_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3278_inst_ack_0, ack => zeropad3D_CP_2067_elements(1048)); -- 
    -- CP-element group 1049:  transition  input  bypass 
    -- CP-element group 1049: predecessors 
    -- CP-element group 1049: 	499 
    -- CP-element group 1049: successors 
    -- CP-element group 1049: 	1050 
    -- CP-element group 1049:  members (2) 
      -- CP-element group 1049: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/Update/$exit
      -- CP-element group 1049: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/Update/ca
      -- 
    ca_12571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1049_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3278_inst_ack_1, ack => zeropad3D_CP_2067_elements(1049)); -- 
    -- CP-element group 1050:  join  transition  output  bypass 
    -- CP-element group 1050: predecessors 
    -- CP-element group 1050: 	1048 
    -- CP-element group 1050: 	1049 
    -- CP-element group 1050: successors 
    -- CP-element group 1050: 	1055 
    -- CP-element group 1050:  members (5) 
      -- CP-element group 1050: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/$exit
      -- CP-element group 1050: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/$exit
      -- CP-element group 1050: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/$exit
      -- CP-element group 1050: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3278/SplitProtocol/$exit
      -- CP-element group 1050: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_req
      -- 
    phi_stmt_3275_req_12572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3275_req_12572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1050), ack => phi_stmt_3275_req_0); -- 
    zeropad3D_cp_element_group_1050: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1050"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1048) & zeropad3D_CP_2067_elements(1049);
      gj_zeropad3D_cp_element_group_1050 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1050), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1051:  transition  input  bypass 
    -- CP-element group 1051: predecessors 
    -- CP-element group 1051: 	499 
    -- CP-element group 1051: successors 
    -- CP-element group 1051: 	1053 
    -- CP-element group 1051:  members (2) 
      -- CP-element group 1051: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/Sample/$exit
      -- CP-element group 1051: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/Sample/ra
      -- 
    ra_12589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1051_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3274_inst_ack_0, ack => zeropad3D_CP_2067_elements(1051)); -- 
    -- CP-element group 1052:  transition  input  bypass 
    -- CP-element group 1052: predecessors 
    -- CP-element group 1052: 	499 
    -- CP-element group 1052: successors 
    -- CP-element group 1052: 	1053 
    -- CP-element group 1052:  members (2) 
      -- CP-element group 1052: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/Update/$exit
      -- CP-element group 1052: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/Update/ca
      -- 
    ca_12594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1052_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3274_inst_ack_1, ack => zeropad3D_CP_2067_elements(1052)); -- 
    -- CP-element group 1053:  join  transition  output  bypass 
    -- CP-element group 1053: predecessors 
    -- CP-element group 1053: 	1051 
    -- CP-element group 1053: 	1052 
    -- CP-element group 1053: successors 
    -- CP-element group 1053: 	1055 
    -- CP-element group 1053:  members (5) 
      -- CP-element group 1053: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/$exit
      -- CP-element group 1053: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/$exit
      -- CP-element group 1053: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/$exit
      -- CP-element group 1053: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3274/SplitProtocol/$exit
      -- CP-element group 1053: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_req
      -- 
    phi_stmt_3269_req_12595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3269_req_12595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1053), ack => phi_stmt_3269_req_1); -- 
    zeropad3D_cp_element_group_1053: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1053"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1051) & zeropad3D_CP_2067_elements(1052);
      gj_zeropad3D_cp_element_group_1053 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1053), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1054:  transition  output  delay-element  bypass 
    -- CP-element group 1054: predecessors 
    -- CP-element group 1054: 	499 
    -- CP-element group 1054: successors 
    -- CP-element group 1054: 	1055 
    -- CP-element group 1054:  members (4) 
      -- CP-element group 1054: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3262/$exit
      -- CP-element group 1054: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/$exit
      -- CP-element group 1054: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3266_konst_delay_trans
      -- CP-element group 1054: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_req
      -- 
    phi_stmt_3262_req_12603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3262_req_12603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1054), ack => phi_stmt_3262_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(1054) is a control-delay.
    cp_element_1054_delay: control_delay_element  generic map(name => " 1054_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(499), ack => zeropad3D_CP_2067_elements(1054), clk => clk, reset =>reset);
    -- CP-element group 1055:  join  transition  bypass 
    -- CP-element group 1055: predecessors 
    -- CP-element group 1055: 	1050 
    -- CP-element group 1055: 	1053 
    -- CP-element group 1055: 	1054 
    -- CP-element group 1055: successors 
    -- CP-element group 1055: 	1066 
    -- CP-element group 1055:  members (1) 
      -- CP-element group 1055: 	 branch_block_stmt_655/ifx_xelse1009_ifx_xend1047_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1055: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1055"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1050) & zeropad3D_CP_2067_elements(1053) & zeropad3D_CP_2067_elements(1054);
      gj_zeropad3D_cp_element_group_1055 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1055), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1056:  transition  input  bypass 
    -- CP-element group 1056: predecessors 
    -- CP-element group 1056: 	480 
    -- CP-element group 1056: successors 
    -- CP-element group 1056: 	1058 
    -- CP-element group 1056:  members (2) 
      -- CP-element group 1056: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/Sample/$exit
      -- CP-element group 1056: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/Sample/ra
      -- 
    ra_12623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1056_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3280_inst_ack_0, ack => zeropad3D_CP_2067_elements(1056)); -- 
    -- CP-element group 1057:  transition  input  bypass 
    -- CP-element group 1057: predecessors 
    -- CP-element group 1057: 	480 
    -- CP-element group 1057: successors 
    -- CP-element group 1057: 	1058 
    -- CP-element group 1057:  members (2) 
      -- CP-element group 1057: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/Update/$exit
      -- CP-element group 1057: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/Update/ca
      -- 
    ca_12628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1057_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3280_inst_ack_1, ack => zeropad3D_CP_2067_elements(1057)); -- 
    -- CP-element group 1058:  join  transition  output  bypass 
    -- CP-element group 1058: predecessors 
    -- CP-element group 1058: 	1056 
    -- CP-element group 1058: 	1057 
    -- CP-element group 1058: successors 
    -- CP-element group 1058: 	1065 
    -- CP-element group 1058:  members (5) 
      -- CP-element group 1058: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/$exit
      -- CP-element group 1058: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/$exit
      -- CP-element group 1058: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/$exit
      -- CP-element group 1058: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_sources/type_cast_3280/SplitProtocol/$exit
      -- CP-element group 1058: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3275/phi_stmt_3275_req
      -- 
    phi_stmt_3275_req_12629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3275_req_12629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1058), ack => phi_stmt_3275_req_1); -- 
    zeropad3D_cp_element_group_1058: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1058"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1056) & zeropad3D_CP_2067_elements(1057);
      gj_zeropad3D_cp_element_group_1058 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1058), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1059:  transition  input  bypass 
    -- CP-element group 1059: predecessors 
    -- CP-element group 1059: 	480 
    -- CP-element group 1059: successors 
    -- CP-element group 1059: 	1061 
    -- CP-element group 1059:  members (2) 
      -- CP-element group 1059: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/Sample/$exit
      -- CP-element group 1059: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/Sample/ra
      -- 
    ra_12646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1059_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3272_inst_ack_0, ack => zeropad3D_CP_2067_elements(1059)); -- 
    -- CP-element group 1060:  transition  input  bypass 
    -- CP-element group 1060: predecessors 
    -- CP-element group 1060: 	480 
    -- CP-element group 1060: successors 
    -- CP-element group 1060: 	1061 
    -- CP-element group 1060:  members (2) 
      -- CP-element group 1060: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/Update/$exit
      -- CP-element group 1060: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/Update/ca
      -- 
    ca_12651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1060_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3272_inst_ack_1, ack => zeropad3D_CP_2067_elements(1060)); -- 
    -- CP-element group 1061:  join  transition  output  bypass 
    -- CP-element group 1061: predecessors 
    -- CP-element group 1061: 	1059 
    -- CP-element group 1061: 	1060 
    -- CP-element group 1061: successors 
    -- CP-element group 1061: 	1065 
    -- CP-element group 1061:  members (5) 
      -- CP-element group 1061: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/$exit
      -- CP-element group 1061: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/$exit
      -- CP-element group 1061: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/$exit
      -- CP-element group 1061: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_sources/type_cast_3272/SplitProtocol/$exit
      -- CP-element group 1061: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3269/phi_stmt_3269_req
      -- 
    phi_stmt_3269_req_12652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3269_req_12652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1061), ack => phi_stmt_3269_req_0); -- 
    zeropad3D_cp_element_group_1061: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1061"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1059) & zeropad3D_CP_2067_elements(1060);
      gj_zeropad3D_cp_element_group_1061 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1061), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1062:  transition  input  bypass 
    -- CP-element group 1062: predecessors 
    -- CP-element group 1062: 	480 
    -- CP-element group 1062: successors 
    -- CP-element group 1062: 	1064 
    -- CP-element group 1062:  members (2) 
      -- CP-element group 1062: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/Sample/$exit
      -- CP-element group 1062: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/Sample/ra
      -- 
    ra_12669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1062_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3268_inst_ack_0, ack => zeropad3D_CP_2067_elements(1062)); -- 
    -- CP-element group 1063:  transition  input  bypass 
    -- CP-element group 1063: predecessors 
    -- CP-element group 1063: 	480 
    -- CP-element group 1063: successors 
    -- CP-element group 1063: 	1064 
    -- CP-element group 1063:  members (2) 
      -- CP-element group 1063: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/Update/$exit
      -- CP-element group 1063: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/Update/ca
      -- 
    ca_12674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1063_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3268_inst_ack_1, ack => zeropad3D_CP_2067_elements(1063)); -- 
    -- CP-element group 1064:  join  transition  output  bypass 
    -- CP-element group 1064: predecessors 
    -- CP-element group 1064: 	1062 
    -- CP-element group 1064: 	1063 
    -- CP-element group 1064: successors 
    -- CP-element group 1064: 	1065 
    -- CP-element group 1064:  members (5) 
      -- CP-element group 1064: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/$exit
      -- CP-element group 1064: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/$exit
      -- CP-element group 1064: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/$exit
      -- CP-element group 1064: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_sources/type_cast_3268/SplitProtocol/$exit
      -- CP-element group 1064: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/phi_stmt_3262/phi_stmt_3262_req
      -- 
    phi_stmt_3262_req_12675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3262_req_12675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1064), ack => phi_stmt_3262_req_1); -- 
    zeropad3D_cp_element_group_1064: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1064"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1062) & zeropad3D_CP_2067_elements(1063);
      gj_zeropad3D_cp_element_group_1064 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1064), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1065:  join  transition  bypass 
    -- CP-element group 1065: predecessors 
    -- CP-element group 1065: 	1058 
    -- CP-element group 1065: 	1061 
    -- CP-element group 1065: 	1064 
    -- CP-element group 1065: successors 
    -- CP-element group 1065: 	1066 
    -- CP-element group 1065:  members (1) 
      -- CP-element group 1065: 	 branch_block_stmt_655/ifx_xthen1004_ifx_xend1047_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1065: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1065"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1058) & zeropad3D_CP_2067_elements(1061) & zeropad3D_CP_2067_elements(1064);
      gj_zeropad3D_cp_element_group_1065 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1065), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1066:  merge  fork  transition  place  bypass 
    -- CP-element group 1066: predecessors 
    -- CP-element group 1066: 	1055 
    -- CP-element group 1066: 	1065 
    -- CP-element group 1066: successors 
    -- CP-element group 1066: 	1067 
    -- CP-element group 1066: 	1068 
    -- CP-element group 1066: 	1069 
    -- CP-element group 1066:  members (2) 
      -- CP-element group 1066: 	 branch_block_stmt_655/merge_stmt_3261_PhiReqMerge
      -- CP-element group 1066: 	 branch_block_stmt_655/merge_stmt_3261_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1066) <= OrReduce(zeropad3D_CP_2067_elements(1055) & zeropad3D_CP_2067_elements(1065));
    -- CP-element group 1067:  transition  input  bypass 
    -- CP-element group 1067: predecessors 
    -- CP-element group 1067: 	1066 
    -- CP-element group 1067: successors 
    -- CP-element group 1067: 	1070 
    -- CP-element group 1067:  members (1) 
      -- CP-element group 1067: 	 branch_block_stmt_655/merge_stmt_3261_PhiAck/phi_stmt_3262_ack
      -- 
    phi_stmt_3262_ack_12680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1067_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3262_ack_0, ack => zeropad3D_CP_2067_elements(1067)); -- 
    -- CP-element group 1068:  transition  input  bypass 
    -- CP-element group 1068: predecessors 
    -- CP-element group 1068: 	1066 
    -- CP-element group 1068: successors 
    -- CP-element group 1068: 	1070 
    -- CP-element group 1068:  members (1) 
      -- CP-element group 1068: 	 branch_block_stmt_655/merge_stmt_3261_PhiAck/phi_stmt_3269_ack
      -- 
    phi_stmt_3269_ack_12681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1068_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3269_ack_0, ack => zeropad3D_CP_2067_elements(1068)); -- 
    -- CP-element group 1069:  transition  input  bypass 
    -- CP-element group 1069: predecessors 
    -- CP-element group 1069: 	1066 
    -- CP-element group 1069: successors 
    -- CP-element group 1069: 	1070 
    -- CP-element group 1069:  members (1) 
      -- CP-element group 1069: 	 branch_block_stmt_655/merge_stmt_3261_PhiAck/phi_stmt_3275_ack
      -- 
    phi_stmt_3275_ack_12682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1069_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3275_ack_0, ack => zeropad3D_CP_2067_elements(1069)); -- 
    -- CP-element group 1070:  join  transition  bypass 
    -- CP-element group 1070: predecessors 
    -- CP-element group 1070: 	1067 
    -- CP-element group 1070: 	1068 
    -- CP-element group 1070: 	1069 
    -- CP-element group 1070: successors 
    -- CP-element group 1070: 	5 
    -- CP-element group 1070:  members (1) 
      -- CP-element group 1070: 	 branch_block_stmt_655/merge_stmt_3261_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1070: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1070"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1067) & zeropad3D_CP_2067_elements(1068) & zeropad3D_CP_2067_elements(1069);
      gj_zeropad3D_cp_element_group_1070 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1070), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1071:  transition  input  bypass 
    -- CP-element group 1071: predecessors 
    -- CP-element group 1071: 	498 
    -- CP-element group 1071: successors 
    -- CP-element group 1071: 	1073 
    -- CP-element group 1071:  members (2) 
      -- CP-element group 1071: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/Sample/$exit
      -- CP-element group 1071: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/Sample/ra
      -- 
    ra_12702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1071_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3295_inst_ack_0, ack => zeropad3D_CP_2067_elements(1071)); -- 
    -- CP-element group 1072:  transition  input  bypass 
    -- CP-element group 1072: predecessors 
    -- CP-element group 1072: 	498 
    -- CP-element group 1072: successors 
    -- CP-element group 1072: 	1073 
    -- CP-element group 1072:  members (2) 
      -- CP-element group 1072: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/Update/$exit
      -- CP-element group 1072: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/Update/ca
      -- 
    ca_12707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1072_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3295_inst_ack_1, ack => zeropad3D_CP_2067_elements(1072)); -- 
    -- CP-element group 1073:  join  transition  output  bypass 
    -- CP-element group 1073: predecessors 
    -- CP-element group 1073: 	1071 
    -- CP-element group 1073: 	1072 
    -- CP-element group 1073: successors 
    -- CP-element group 1073: 	1080 
    -- CP-element group 1073:  members (5) 
      -- CP-element group 1073: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/$exit
      -- CP-element group 1073: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/$exit
      -- CP-element group 1073: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/$exit
      -- CP-element group 1073: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_sources/type_cast_3295/SplitProtocol/$exit
      -- CP-element group 1073: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3292/phi_stmt_3292_req
      -- 
    phi_stmt_3292_req_12708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3292_req_12708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1073), ack => phi_stmt_3292_req_0); -- 
    zeropad3D_cp_element_group_1073: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1073"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1071) & zeropad3D_CP_2067_elements(1072);
      gj_zeropad3D_cp_element_group_1073 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1073), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1074:  transition  input  bypass 
    -- CP-element group 1074: predecessors 
    -- CP-element group 1074: 	498 
    -- CP-element group 1074: successors 
    -- CP-element group 1074: 	1076 
    -- CP-element group 1074:  members (2) 
      -- CP-element group 1074: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/Sample/$exit
      -- CP-element group 1074: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/Sample/ra
      -- 
    ra_12725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1074_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3291_inst_ack_0, ack => zeropad3D_CP_2067_elements(1074)); -- 
    -- CP-element group 1075:  transition  input  bypass 
    -- CP-element group 1075: predecessors 
    -- CP-element group 1075: 	498 
    -- CP-element group 1075: successors 
    -- CP-element group 1075: 	1076 
    -- CP-element group 1075:  members (2) 
      -- CP-element group 1075: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/Update/$exit
      -- CP-element group 1075: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/Update/ca
      -- 
    ca_12730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1075_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3291_inst_ack_1, ack => zeropad3D_CP_2067_elements(1075)); -- 
    -- CP-element group 1076:  join  transition  output  bypass 
    -- CP-element group 1076: predecessors 
    -- CP-element group 1076: 	1074 
    -- CP-element group 1076: 	1075 
    -- CP-element group 1076: successors 
    -- CP-element group 1076: 	1080 
    -- CP-element group 1076:  members (5) 
      -- CP-element group 1076: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/$exit
      -- CP-element group 1076: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/$exit
      -- CP-element group 1076: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/$exit
      -- CP-element group 1076: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_sources/type_cast_3291/SplitProtocol/$exit
      -- CP-element group 1076: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3288/phi_stmt_3288_req
      -- 
    phi_stmt_3288_req_12731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3288_req_12731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1076), ack => phi_stmt_3288_req_0); -- 
    zeropad3D_cp_element_group_1076: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1076"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1074) & zeropad3D_CP_2067_elements(1075);
      gj_zeropad3D_cp_element_group_1076 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1076), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1077:  transition  input  bypass 
    -- CP-element group 1077: predecessors 
    -- CP-element group 1077: 	498 
    -- CP-element group 1077: successors 
    -- CP-element group 1077: 	1079 
    -- CP-element group 1077:  members (2) 
      -- CP-element group 1077: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/Sample/$exit
      -- CP-element group 1077: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/Sample/ra
      -- 
    ra_12748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1077_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3287_inst_ack_0, ack => zeropad3D_CP_2067_elements(1077)); -- 
    -- CP-element group 1078:  transition  input  bypass 
    -- CP-element group 1078: predecessors 
    -- CP-element group 1078: 	498 
    -- CP-element group 1078: successors 
    -- CP-element group 1078: 	1079 
    -- CP-element group 1078:  members (2) 
      -- CP-element group 1078: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/Update/$exit
      -- CP-element group 1078: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/Update/ca
      -- 
    ca_12753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1078_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3287_inst_ack_1, ack => zeropad3D_CP_2067_elements(1078)); -- 
    -- CP-element group 1079:  join  transition  output  bypass 
    -- CP-element group 1079: predecessors 
    -- CP-element group 1079: 	1077 
    -- CP-element group 1079: 	1078 
    -- CP-element group 1079: successors 
    -- CP-element group 1079: 	1080 
    -- CP-element group 1079:  members (5) 
      -- CP-element group 1079: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/$exit
      -- CP-element group 1079: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/$exit
      -- CP-element group 1079: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/$exit
      -- CP-element group 1079: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_sources/type_cast_3287/SplitProtocol/$exit
      -- CP-element group 1079: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/phi_stmt_3284/phi_stmt_3284_req
      -- 
    phi_stmt_3284_req_12754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3284_req_12754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1079), ack => phi_stmt_3284_req_0); -- 
    zeropad3D_cp_element_group_1079: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1079"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1077) & zeropad3D_CP_2067_elements(1078);
      gj_zeropad3D_cp_element_group_1079 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1079), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1080:  join  fork  transition  place  bypass 
    -- CP-element group 1080: predecessors 
    -- CP-element group 1080: 	1073 
    -- CP-element group 1080: 	1076 
    -- CP-element group 1080: 	1079 
    -- CP-element group 1080: successors 
    -- CP-element group 1080: 	1081 
    -- CP-element group 1080: 	1082 
    -- CP-element group 1080: 	1083 
    -- CP-element group 1080:  members (3) 
      -- CP-element group 1080: 	 branch_block_stmt_655/ifx_xelse1009_whilex_xend1048_PhiReq/$exit
      -- CP-element group 1080: 	 branch_block_stmt_655/merge_stmt_3283_PhiReqMerge
      -- CP-element group 1080: 	 branch_block_stmt_655/merge_stmt_3283_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_1080: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1080"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1073) & zeropad3D_CP_2067_elements(1076) & zeropad3D_CP_2067_elements(1079);
      gj_zeropad3D_cp_element_group_1080 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1080), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1081:  transition  input  bypass 
    -- CP-element group 1081: predecessors 
    -- CP-element group 1081: 	1080 
    -- CP-element group 1081: successors 
    -- CP-element group 1081: 	1084 
    -- CP-element group 1081:  members (1) 
      -- CP-element group 1081: 	 branch_block_stmt_655/merge_stmt_3283_PhiAck/phi_stmt_3284_ack
      -- 
    phi_stmt_3284_ack_12759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1081_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3284_ack_0, ack => zeropad3D_CP_2067_elements(1081)); -- 
    -- CP-element group 1082:  transition  input  bypass 
    -- CP-element group 1082: predecessors 
    -- CP-element group 1082: 	1080 
    -- CP-element group 1082: successors 
    -- CP-element group 1082: 	1084 
    -- CP-element group 1082:  members (1) 
      -- CP-element group 1082: 	 branch_block_stmt_655/merge_stmt_3283_PhiAck/phi_stmt_3288_ack
      -- 
    phi_stmt_3288_ack_12760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1082_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3288_ack_0, ack => zeropad3D_CP_2067_elements(1082)); -- 
    -- CP-element group 1083:  transition  input  bypass 
    -- CP-element group 1083: predecessors 
    -- CP-element group 1083: 	1080 
    -- CP-element group 1083: successors 
    -- CP-element group 1083: 	1084 
    -- CP-element group 1083:  members (1) 
      -- CP-element group 1083: 	 branch_block_stmt_655/merge_stmt_3283_PhiAck/phi_stmt_3292_ack
      -- 
    phi_stmt_3292_ack_12761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1083_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3292_ack_0, ack => zeropad3D_CP_2067_elements(1083)); -- 
    -- CP-element group 1084:  join  fork  transition  place  output  bypass 
    -- CP-element group 1084: predecessors 
    -- CP-element group 1084: 	1081 
    -- CP-element group 1084: 	1082 
    -- CP-element group 1084: 	1083 
    -- CP-element group 1084: successors 
    -- CP-element group 1084: 	500 
    -- CP-element group 1084: 	501 
    -- CP-element group 1084: 	502 
    -- CP-element group 1084: 	503 
    -- CP-element group 1084: 	504 
    -- CP-element group 1084: 	505 
    -- CP-element group 1084: 	506 
    -- CP-element group 1084: 	507 
    -- CP-element group 1084: 	508 
    -- CP-element group 1084: 	509 
    -- CP-element group 1084: 	510 
    -- CP-element group 1084: 	511 
    -- CP-element group 1084: 	513 
    -- CP-element group 1084: 	515 
    -- CP-element group 1084: 	517 
    -- CP-element group 1084: 	519 
    -- CP-element group 1084: 	521 
    -- CP-element group 1084:  members (79) 
      -- CP-element group 1084: 	 branch_block_stmt_655/merge_stmt_3283__exit__
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394__entry__
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_Update/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_Update/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3339_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_Update/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3335_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3352_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_Update/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_Update/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3348_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_sample_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_Sample/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_Sample/rr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3299_Update/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_sample_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_Sample/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_Sample/rr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3309_Update/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_sample_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_word_address_calculated
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_root_address_calculated
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Sample/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Sample/word_access_start/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Sample/word_access_start/word_0/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Sample/word_access_start/word_0/rr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/word_access_complete/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/word_access_complete/word_0/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_pad_3318_Update/word_access_complete/word_0/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_sample_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_word_address_calculated
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_root_address_calculated
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Sample/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Sample/word_access_start/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Sample/word_access_start/word_0/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Sample/word_access_start/word_0/rr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/word_access_complete/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/word_access_complete/word_0/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_depth_high_3321_Update/word_access_complete/word_0/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_sample_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_word_address_calculated
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_root_address_calculated
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Sample/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Sample/word_access_start/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Sample/word_access_start/word_0/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Sample/word_access_start/word_0/rr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/word_access_complete/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/word_access_complete/word_0/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_depth_high_3324_Update/word_access_complete/word_0/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_sample_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_word_address_calculated
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_root_address_calculated
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Sample/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Sample/word_access_start/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Sample/word_access_start/word_0/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Sample/word_access_start/word_0/rr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/word_access_complete/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/word_access_complete/word_0/$entry
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/LOAD_out_col_high_3327_Update/word_access_complete/word_0/cr
      -- CP-element group 1084: 	 branch_block_stmt_655/assign_stmt_3300_to_assign_stmt_3394/type_cast_3331_update_start_
      -- CP-element group 1084: 	 branch_block_stmt_655/merge_stmt_3283_PhiAck/$exit
      -- 
    cr_7828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3352_inst_req_1); -- 
    cr_7800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3339_inst_req_1); -- 
    cr_7786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3335_inst_req_1); -- 
    cr_7772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3331_inst_req_1); -- 
    cr_7814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3348_inst_req_1); -- 
    rr_7607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3299_inst_req_0); -- 
    cr_7612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3299_inst_req_1); -- 
    rr_7621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3309_inst_req_0); -- 
    cr_7626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => type_cast_3309_inst_req_1); -- 
    rr_7643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => LOAD_pad_3318_load_0_req_0); -- 
    cr_7654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => LOAD_pad_3318_load_0_req_1); -- 
    rr_7676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => LOAD_depth_high_3321_load_0_req_0); -- 
    cr_7687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => LOAD_depth_high_3321_load_0_req_1); -- 
    rr_7709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => LOAD_out_depth_high_3324_load_0_req_0); -- 
    cr_7720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => LOAD_out_depth_high_3324_load_0_req_1); -- 
    rr_7742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => LOAD_out_col_high_3327_load_0_req_0); -- 
    cr_7753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1084), ack => LOAD_out_col_high_3327_load_0_req_1); -- 
    zeropad3D_cp_element_group_1084: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1084"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1081) & zeropad3D_CP_2067_elements(1082) & zeropad3D_CP_2067_elements(1083);
      gj_zeropad3D_cp_element_group_1084 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1084), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1085:  transition  input  bypass 
    -- CP-element group 1085: predecessors 
    -- CP-element group 1085: 	6 
    -- CP-element group 1085: successors 
    -- CP-element group 1085: 	1087 
    -- CP-element group 1085:  members (2) 
      -- CP-element group 1085: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/Sample/$exit
      -- CP-element group 1085: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/Sample/ra
      -- 
    ra_12781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1085_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3403_inst_ack_0, ack => zeropad3D_CP_2067_elements(1085)); -- 
    -- CP-element group 1086:  transition  input  bypass 
    -- CP-element group 1086: predecessors 
    -- CP-element group 1086: 	6 
    -- CP-element group 1086: successors 
    -- CP-element group 1086: 	1087 
    -- CP-element group 1086:  members (2) 
      -- CP-element group 1086: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/Update/$exit
      -- CP-element group 1086: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/Update/ca
      -- 
    ca_12786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1086_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3403_inst_ack_1, ack => zeropad3D_CP_2067_elements(1086)); -- 
    -- CP-element group 1087:  join  transition  output  bypass 
    -- CP-element group 1087: predecessors 
    -- CP-element group 1087: 	1085 
    -- CP-element group 1087: 	1086 
    -- CP-element group 1087: successors 
    -- CP-element group 1087: 	1094 
    -- CP-element group 1087:  members (5) 
      -- CP-element group 1087: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/$exit
      -- CP-element group 1087: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/$exit
      -- CP-element group 1087: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/$exit
      -- CP-element group 1087: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3403/SplitProtocol/$exit
      -- CP-element group 1087: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_req
      -- 
    phi_stmt_3397_req_12787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3397_req_12787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1087), ack => phi_stmt_3397_req_1); -- 
    zeropad3D_cp_element_group_1087: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1087"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1085) & zeropad3D_CP_2067_elements(1086);
      gj_zeropad3D_cp_element_group_1087 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1087), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1088:  transition  input  bypass 
    -- CP-element group 1088: predecessors 
    -- CP-element group 1088: 	6 
    -- CP-element group 1088: successors 
    -- CP-element group 1088: 	1090 
    -- CP-element group 1088:  members (2) 
      -- CP-element group 1088: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/Sample/$exit
      -- CP-element group 1088: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/Sample/ra
      -- 
    ra_12804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1088_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3407_inst_ack_0, ack => zeropad3D_CP_2067_elements(1088)); -- 
    -- CP-element group 1089:  transition  input  bypass 
    -- CP-element group 1089: predecessors 
    -- CP-element group 1089: 	6 
    -- CP-element group 1089: successors 
    -- CP-element group 1089: 	1090 
    -- CP-element group 1089:  members (2) 
      -- CP-element group 1089: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/Update/ca
      -- CP-element group 1089: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/Update/$exit
      -- 
    ca_12809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1089_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3407_inst_ack_1, ack => zeropad3D_CP_2067_elements(1089)); -- 
    -- CP-element group 1090:  join  transition  output  bypass 
    -- CP-element group 1090: predecessors 
    -- CP-element group 1090: 	1088 
    -- CP-element group 1090: 	1089 
    -- CP-element group 1090: successors 
    -- CP-element group 1090: 	1094 
    -- CP-element group 1090:  members (5) 
      -- CP-element group 1090: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_req
      -- CP-element group 1090: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/$exit
      -- CP-element group 1090: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/$exit
      -- CP-element group 1090: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/$exit
      -- CP-element group 1090: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3407/SplitProtocol/$exit
      -- 
    phi_stmt_3404_req_12810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3404_req_12810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1090), ack => phi_stmt_3404_req_0); -- 
    zeropad3D_cp_element_group_1090: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1090"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1088) & zeropad3D_CP_2067_elements(1089);
      gj_zeropad3D_cp_element_group_1090 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1090), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1091:  transition  input  bypass 
    -- CP-element group 1091: predecessors 
    -- CP-element group 1091: 	6 
    -- CP-element group 1091: successors 
    -- CP-element group 1091: 	1093 
    -- CP-element group 1091:  members (2) 
      -- CP-element group 1091: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/Sample/ra
      -- CP-element group 1091: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/Sample/$exit
      -- 
    ra_12827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1091_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3415_inst_ack_0, ack => zeropad3D_CP_2067_elements(1091)); -- 
    -- CP-element group 1092:  transition  input  bypass 
    -- CP-element group 1092: predecessors 
    -- CP-element group 1092: 	6 
    -- CP-element group 1092: successors 
    -- CP-element group 1092: 	1093 
    -- CP-element group 1092:  members (2) 
      -- CP-element group 1092: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/Update/ca
      -- CP-element group 1092: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/Update/$exit
      -- 
    ca_12832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1092_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3415_inst_ack_1, ack => zeropad3D_CP_2067_elements(1092)); -- 
    -- CP-element group 1093:  join  transition  output  bypass 
    -- CP-element group 1093: predecessors 
    -- CP-element group 1093: 	1091 
    -- CP-element group 1093: 	1092 
    -- CP-element group 1093: successors 
    -- CP-element group 1093: 	1094 
    -- CP-element group 1093:  members (5) 
      -- CP-element group 1093: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/$exit
      -- CP-element group 1093: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_req
      -- CP-element group 1093: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/$exit
      -- CP-element group 1093: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/SplitProtocol/$exit
      -- CP-element group 1093: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3415/$exit
      -- 
    phi_stmt_3410_req_12833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3410_req_12833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1093), ack => phi_stmt_3410_req_1); -- 
    zeropad3D_cp_element_group_1093: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1093"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1091) & zeropad3D_CP_2067_elements(1092);
      gj_zeropad3D_cp_element_group_1093 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1093), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1094:  join  transition  bypass 
    -- CP-element group 1094: predecessors 
    -- CP-element group 1094: 	1087 
    -- CP-element group 1094: 	1090 
    -- CP-element group 1094: 	1093 
    -- CP-element group 1094: successors 
    -- CP-element group 1094: 	1103 
    -- CP-element group 1094:  members (1) 
      -- CP-element group 1094: 	 branch_block_stmt_655/ifx_xend1269_whilex_xbody1112_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1094: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1094"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1087) & zeropad3D_CP_2067_elements(1090) & zeropad3D_CP_2067_elements(1093);
      gj_zeropad3D_cp_element_group_1094 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1094), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1095:  transition  output  delay-element  bypass 
    -- CP-element group 1095: predecessors 
    -- CP-element group 1095: 	522 
    -- CP-element group 1095: successors 
    -- CP-element group 1095: 	1102 
    -- CP-element group 1095:  members (4) 
      -- CP-element group 1095: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_req
      -- CP-element group 1095: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/type_cast_3401_konst_delay_trans
      -- CP-element group 1095: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3397/phi_stmt_3397_sources/$exit
      -- CP-element group 1095: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3397/$exit
      -- 
    phi_stmt_3397_req_12844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3397_req_12844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1095), ack => phi_stmt_3397_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(1095) is a control-delay.
    cp_element_1095_delay: control_delay_element  generic map(name => " 1095_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(522), ack => zeropad3D_CP_2067_elements(1095), clk => clk, reset =>reset);
    -- CP-element group 1096:  transition  input  bypass 
    -- CP-element group 1096: predecessors 
    -- CP-element group 1096: 	522 
    -- CP-element group 1096: successors 
    -- CP-element group 1096: 	1098 
    -- CP-element group 1096:  members (2) 
      -- CP-element group 1096: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/Sample/ra
      -- CP-element group 1096: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/Sample/$exit
      -- 
    ra_12861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1096_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3409_inst_ack_0, ack => zeropad3D_CP_2067_elements(1096)); -- 
    -- CP-element group 1097:  transition  input  bypass 
    -- CP-element group 1097: predecessors 
    -- CP-element group 1097: 	522 
    -- CP-element group 1097: successors 
    -- CP-element group 1097: 	1098 
    -- CP-element group 1097:  members (2) 
      -- CP-element group 1097: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/Update/$exit
      -- CP-element group 1097: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/Update/ca
      -- 
    ca_12866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1097_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3409_inst_ack_1, ack => zeropad3D_CP_2067_elements(1097)); -- 
    -- CP-element group 1098:  join  transition  output  bypass 
    -- CP-element group 1098: predecessors 
    -- CP-element group 1098: 	1096 
    -- CP-element group 1098: 	1097 
    -- CP-element group 1098: successors 
    -- CP-element group 1098: 	1102 
    -- CP-element group 1098:  members (5) 
      -- CP-element group 1098: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/SplitProtocol/$exit
      -- CP-element group 1098: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/type_cast_3409/$exit
      -- CP-element group 1098: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_sources/$exit
      -- CP-element group 1098: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/$exit
      -- CP-element group 1098: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3404/phi_stmt_3404_req
      -- 
    phi_stmt_3404_req_12867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3404_req_12867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1098), ack => phi_stmt_3404_req_1); -- 
    zeropad3D_cp_element_group_1098: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1098"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1096) & zeropad3D_CP_2067_elements(1097);
      gj_zeropad3D_cp_element_group_1098 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1098), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1099:  transition  input  bypass 
    -- CP-element group 1099: predecessors 
    -- CP-element group 1099: 	522 
    -- CP-element group 1099: successors 
    -- CP-element group 1099: 	1101 
    -- CP-element group 1099:  members (2) 
      -- CP-element group 1099: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/Sample/ra
      -- CP-element group 1099: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/Sample/$exit
      -- 
    ra_12884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1099_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3413_inst_ack_0, ack => zeropad3D_CP_2067_elements(1099)); -- 
    -- CP-element group 1100:  transition  input  bypass 
    -- CP-element group 1100: predecessors 
    -- CP-element group 1100: 	522 
    -- CP-element group 1100: successors 
    -- CP-element group 1100: 	1101 
    -- CP-element group 1100:  members (2) 
      -- CP-element group 1100: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/Update/$exit
      -- CP-element group 1100: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/Update/ca
      -- 
    ca_12889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3413_inst_ack_1, ack => zeropad3D_CP_2067_elements(1100)); -- 
    -- CP-element group 1101:  join  transition  output  bypass 
    -- CP-element group 1101: predecessors 
    -- CP-element group 1101: 	1099 
    -- CP-element group 1101: 	1100 
    -- CP-element group 1101: successors 
    -- CP-element group 1101: 	1102 
    -- CP-element group 1101:  members (5) 
      -- CP-element group 1101: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/SplitProtocol/$exit
      -- CP-element group 1101: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/type_cast_3413/$exit
      -- CP-element group 1101: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_sources/$exit
      -- CP-element group 1101: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/$exit
      -- CP-element group 1101: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/phi_stmt_3410/phi_stmt_3410_req
      -- 
    phi_stmt_3410_req_12890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3410_req_12890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1101), ack => phi_stmt_3410_req_0); -- 
    zeropad3D_cp_element_group_1101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1099) & zeropad3D_CP_2067_elements(1100);
      gj_zeropad3D_cp_element_group_1101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1102:  join  transition  bypass 
    -- CP-element group 1102: predecessors 
    -- CP-element group 1102: 	1095 
    -- CP-element group 1102: 	1098 
    -- CP-element group 1102: 	1101 
    -- CP-element group 1102: successors 
    -- CP-element group 1102: 	1103 
    -- CP-element group 1102:  members (1) 
      -- CP-element group 1102: 	 branch_block_stmt_655/whilex_xend1048_whilex_xbody1112_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1102: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1102"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1095) & zeropad3D_CP_2067_elements(1098) & zeropad3D_CP_2067_elements(1101);
      gj_zeropad3D_cp_element_group_1102 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1103:  merge  fork  transition  place  bypass 
    -- CP-element group 1103: predecessors 
    -- CP-element group 1103: 	1094 
    -- CP-element group 1103: 	1102 
    -- CP-element group 1103: successors 
    -- CP-element group 1103: 	1104 
    -- CP-element group 1103: 	1105 
    -- CP-element group 1103: 	1106 
    -- CP-element group 1103:  members (2) 
      -- CP-element group 1103: 	 branch_block_stmt_655/merge_stmt_3396_PhiReqMerge
      -- CP-element group 1103: 	 branch_block_stmt_655/merge_stmt_3396_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1103) <= OrReduce(zeropad3D_CP_2067_elements(1094) & zeropad3D_CP_2067_elements(1102));
    -- CP-element group 1104:  transition  input  bypass 
    -- CP-element group 1104: predecessors 
    -- CP-element group 1104: 	1103 
    -- CP-element group 1104: successors 
    -- CP-element group 1104: 	1107 
    -- CP-element group 1104:  members (1) 
      -- CP-element group 1104: 	 branch_block_stmt_655/merge_stmt_3396_PhiAck/phi_stmt_3397_ack
      -- 
    phi_stmt_3397_ack_12895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3397_ack_0, ack => zeropad3D_CP_2067_elements(1104)); -- 
    -- CP-element group 1105:  transition  input  bypass 
    -- CP-element group 1105: predecessors 
    -- CP-element group 1105: 	1103 
    -- CP-element group 1105: successors 
    -- CP-element group 1105: 	1107 
    -- CP-element group 1105:  members (1) 
      -- CP-element group 1105: 	 branch_block_stmt_655/merge_stmt_3396_PhiAck/phi_stmt_3404_ack
      -- 
    phi_stmt_3404_ack_12896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3404_ack_0, ack => zeropad3D_CP_2067_elements(1105)); -- 
    -- CP-element group 1106:  transition  input  bypass 
    -- CP-element group 1106: predecessors 
    -- CP-element group 1106: 	1103 
    -- CP-element group 1106: successors 
    -- CP-element group 1106: 	1107 
    -- CP-element group 1106:  members (1) 
      -- CP-element group 1106: 	 branch_block_stmt_655/merge_stmt_3396_PhiAck/phi_stmt_3410_ack
      -- 
    phi_stmt_3410_ack_12897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3410_ack_0, ack => zeropad3D_CP_2067_elements(1106)); -- 
    -- CP-element group 1107:  join  fork  transition  place  output  bypass 
    -- CP-element group 1107: predecessors 
    -- CP-element group 1107: 	1104 
    -- CP-element group 1107: 	1105 
    -- CP-element group 1107: 	1106 
    -- CP-element group 1107: successors 
    -- CP-element group 1107: 	523 
    -- CP-element group 1107: 	524 
    -- CP-element group 1107:  members (10) 
      -- CP-element group 1107: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428__entry__
      -- CP-element group 1107: 	 branch_block_stmt_655/merge_stmt_3396__exit__
      -- CP-element group 1107: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_Update/cr
      -- CP-element group 1107: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_Update/$entry
      -- CP-element group 1107: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_Sample/rr
      -- CP-element group 1107: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_Sample/$entry
      -- CP-element group 1107: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_update_start_
      -- CP-element group 1107: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/type_cast_3420_sample_start_
      -- CP-element group 1107: 	 branch_block_stmt_655/assign_stmt_3421_to_assign_stmt_3428/$entry
      -- CP-element group 1107: 	 branch_block_stmt_655/merge_stmt_3396_PhiAck/$exit
      -- 
    cr_7845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1107), ack => type_cast_3420_inst_req_1); -- 
    rr_7840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1107), ack => type_cast_3420_inst_req_0); -- 
    zeropad3D_cp_element_group_1107: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1107"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1104) & zeropad3D_CP_2067_elements(1105) & zeropad3D_CP_2067_elements(1106);
      gj_zeropad3D_cp_element_group_1107 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1108:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1108: predecessors 
    -- CP-element group 1108: 	525 
    -- CP-element group 1108: 	532 
    -- CP-element group 1108: 	535 
    -- CP-element group 1108: 	542 
    -- CP-element group 1108: successors 
    -- CP-element group 1108: 	543 
    -- CP-element group 1108: 	544 
    -- CP-element group 1108: 	545 
    -- CP-element group 1108: 	546 
    -- CP-element group 1108: 	549 
    -- CP-element group 1108: 	551 
    -- CP-element group 1108: 	553 
    -- CP-element group 1108: 	555 
    -- CP-element group 1108:  members (33) 
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574__entry__
      -- CP-element group 1108: 	 branch_block_stmt_655/merge_stmt_3518__exit__
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_sample_start_
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_Sample/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_Update/req
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_Update/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_update_start_
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_Update/cr
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_update_start_
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_Update/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_complete/req
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/array_obj_ref_3567_final_index_sum_regn_update_start
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/addr_of_3568_complete/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_Update/cr
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_Sample/rr
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_Update/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3522_update_start_
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3561_update_start_
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_Update/cr
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_Update/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_Sample/rr
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_Sample/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_update_start_
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/type_cast_3527_sample_start_
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Update/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Update/word_access_complete/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Update/word_access_complete/word_0/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/assign_stmt_3523_to_assign_stmt_3574/ptr_deref_3571_Update/word_access_complete/word_0/cr
      -- CP-element group 1108: 	 branch_block_stmt_655/merge_stmt_3518_PhiAck/$entry
      -- CP-element group 1108: 	 branch_block_stmt_655/merge_stmt_3518_PhiReqMerge
      -- CP-element group 1108: 	 branch_block_stmt_655/merge_stmt_3518_PhiAck/$exit
      -- CP-element group 1108: 	 branch_block_stmt_655/merge_stmt_3518_PhiAck/dummy
      -- 
    req_8114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1108), ack => array_obj_ref_3567_index_offset_req_1); -- 
    cr_8055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1108), ack => type_cast_3522_inst_req_1); -- 
    req_8129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1108), ack => addr_of_3568_final_reg_req_1); -- 
    cr_8083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1108), ack => type_cast_3561_inst_req_1); -- 
    rr_8050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1108), ack => type_cast_3522_inst_req_0); -- 
    cr_8069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1108), ack => type_cast_3527_inst_req_1); -- 
    rr_8064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1108), ack => type_cast_3527_inst_req_0); -- 
    cr_8179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1108), ack => ptr_deref_3571_store_0_req_1); -- 
    zeropad3D_CP_2067_elements(1108) <= OrReduce(zeropad3D_CP_2067_elements(525) & zeropad3D_CP_2067_elements(532) & zeropad3D_CP_2067_elements(535) & zeropad3D_CP_2067_elements(542));
    -- CP-element group 1109:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1109: predecessors 
    -- CP-element group 1109: 	556 
    -- CP-element group 1109: 	576 
    -- CP-element group 1109: successors 
    -- CP-element group 1109: 	577 
    -- CP-element group 1109: 	578 
    -- CP-element group 1109:  members (13) 
      -- CP-element group 1109: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701__entry__
      -- CP-element group 1109: 	 branch_block_stmt_655/merge_stmt_3683__exit__
      -- CP-element group 1109: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/$entry
      -- CP-element group 1109: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_sample_start_
      -- CP-element group 1109: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_update_start_
      -- CP-element group 1109: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_Sample/$entry
      -- CP-element group 1109: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_Sample/rr
      -- CP-element group 1109: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_Update/$entry
      -- CP-element group 1109: 	 branch_block_stmt_655/assign_stmt_3688_to_assign_stmt_3701/type_cast_3687_Update/cr
      -- CP-element group 1109: 	 branch_block_stmt_655/merge_stmt_3683_PhiAck/dummy
      -- CP-element group 1109: 	 branch_block_stmt_655/merge_stmt_3683_PhiAck/$exit
      -- CP-element group 1109: 	 branch_block_stmt_655/merge_stmt_3683_PhiAck/$entry
      -- CP-element group 1109: 	 branch_block_stmt_655/merge_stmt_3683_PhiReqMerge
      -- 
    rr_8428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1109), ack => type_cast_3687_inst_req_0); -- 
    cr_8433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1109), ack => type_cast_3687_inst_req_1); -- 
    zeropad3D_CP_2067_elements(1109) <= OrReduce(zeropad3D_CP_2067_elements(556) & zeropad3D_CP_2067_elements(576));
    -- CP-element group 1110:  transition  output  delay-element  bypass 
    -- CP-element group 1110: predecessors 
    -- CP-element group 1110: 	598 
    -- CP-element group 1110: successors 
    -- CP-element group 1110: 	1117 
    -- CP-element group 1110:  members (4) 
      -- CP-element group 1110: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3807_konst_delay_trans
      -- CP-element group 1110: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_req
      -- CP-element group 1110: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/$exit
      -- CP-element group 1110: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3801/$exit
      -- 
    phi_stmt_3801_req_13008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3801_req_13008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1110), ack => phi_stmt_3801_req_1); -- 
    -- Element group zeropad3D_CP_2067_elements(1110) is a control-delay.
    cp_element_1110_delay: control_delay_element  generic map(name => " 1110_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(598), ack => zeropad3D_CP_2067_elements(1110), clk => clk, reset =>reset);
    -- CP-element group 1111:  transition  input  bypass 
    -- CP-element group 1111: predecessors 
    -- CP-element group 1111: 	598 
    -- CP-element group 1111: successors 
    -- CP-element group 1111: 	1113 
    -- CP-element group 1111:  members (2) 
      -- CP-element group 1111: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/Sample/$exit
      -- CP-element group 1111: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/Sample/ra
      -- 
    ra_13025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3813_inst_ack_0, ack => zeropad3D_CP_2067_elements(1111)); -- 
    -- CP-element group 1112:  transition  input  bypass 
    -- CP-element group 1112: predecessors 
    -- CP-element group 1112: 	598 
    -- CP-element group 1112: successors 
    -- CP-element group 1112: 	1113 
    -- CP-element group 1112:  members (2) 
      -- CP-element group 1112: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/Update/ca
      -- CP-element group 1112: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/Update/$exit
      -- 
    ca_13030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3813_inst_ack_1, ack => zeropad3D_CP_2067_elements(1112)); -- 
    -- CP-element group 1113:  join  transition  output  bypass 
    -- CP-element group 1113: predecessors 
    -- CP-element group 1113: 	1111 
    -- CP-element group 1113: 	1112 
    -- CP-element group 1113: successors 
    -- CP-element group 1113: 	1117 
    -- CP-element group 1113:  members (5) 
      -- CP-element group 1113: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_req
      -- CP-element group 1113: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/$exit
      -- CP-element group 1113: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/$exit
      -- CP-element group 1113: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/$exit
      -- CP-element group 1113: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3813/SplitProtocol/$exit
      -- 
    phi_stmt_3808_req_13031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3808_req_13031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1113), ack => phi_stmt_3808_req_1); -- 
    zeropad3D_cp_element_group_1113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1111) & zeropad3D_CP_2067_elements(1112);
      gj_zeropad3D_cp_element_group_1113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1114:  transition  input  bypass 
    -- CP-element group 1114: predecessors 
    -- CP-element group 1114: 	598 
    -- CP-element group 1114: successors 
    -- CP-element group 1114: 	1116 
    -- CP-element group 1114:  members (2) 
      -- CP-element group 1114: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/Sample/ra
      -- CP-element group 1114: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/Sample/$exit
      -- 
    ra_13048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3819_inst_ack_0, ack => zeropad3D_CP_2067_elements(1114)); -- 
    -- CP-element group 1115:  transition  input  bypass 
    -- CP-element group 1115: predecessors 
    -- CP-element group 1115: 	598 
    -- CP-element group 1115: successors 
    -- CP-element group 1115: 	1116 
    -- CP-element group 1115:  members (2) 
      -- CP-element group 1115: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/Update/ca
      -- CP-element group 1115: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/Update/$exit
      -- 
    ca_13053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3819_inst_ack_1, ack => zeropad3D_CP_2067_elements(1115)); -- 
    -- CP-element group 1116:  join  transition  output  bypass 
    -- CP-element group 1116: predecessors 
    -- CP-element group 1116: 	1114 
    -- CP-element group 1116: 	1115 
    -- CP-element group 1116: successors 
    -- CP-element group 1116: 	1117 
    -- CP-element group 1116:  members (5) 
      -- CP-element group 1116: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_req
      -- CP-element group 1116: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/SplitProtocol/$exit
      -- CP-element group 1116: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3819/$exit
      -- CP-element group 1116: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/$exit
      -- CP-element group 1116: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/phi_stmt_3814/$exit
      -- 
    phi_stmt_3814_req_13054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3814_req_13054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1116), ack => phi_stmt_3814_req_1); -- 
    zeropad3D_cp_element_group_1116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1114) & zeropad3D_CP_2067_elements(1115);
      gj_zeropad3D_cp_element_group_1116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1117:  join  transition  bypass 
    -- CP-element group 1117: predecessors 
    -- CP-element group 1117: 	1110 
    -- CP-element group 1117: 	1113 
    -- CP-element group 1117: 	1116 
    -- CP-element group 1117: successors 
    -- CP-element group 1117: 	1128 
    -- CP-element group 1117:  members (1) 
      -- CP-element group 1117: 	 branch_block_stmt_655/ifx_xelse1232_ifx_xend1269_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1110) & zeropad3D_CP_2067_elements(1113) & zeropad3D_CP_2067_elements(1116);
      gj_zeropad3D_cp_element_group_1117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1118:  transition  input  bypass 
    -- CP-element group 1118: predecessors 
    -- CP-element group 1118: 	579 
    -- CP-element group 1118: successors 
    -- CP-element group 1118: 	1120 
    -- CP-element group 1118:  members (2) 
      -- CP-element group 1118: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/Sample/ra
      -- CP-element group 1118: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/Sample/$exit
      -- 
    ra_13074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3804_inst_ack_0, ack => zeropad3D_CP_2067_elements(1118)); -- 
    -- CP-element group 1119:  transition  input  bypass 
    -- CP-element group 1119: predecessors 
    -- CP-element group 1119: 	579 
    -- CP-element group 1119: successors 
    -- CP-element group 1119: 	1120 
    -- CP-element group 1119:  members (2) 
      -- CP-element group 1119: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/Update/$exit
      -- CP-element group 1119: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/Update/ca
      -- 
    ca_13079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3804_inst_ack_1, ack => zeropad3D_CP_2067_elements(1119)); -- 
    -- CP-element group 1120:  join  transition  output  bypass 
    -- CP-element group 1120: predecessors 
    -- CP-element group 1120: 	1118 
    -- CP-element group 1120: 	1119 
    -- CP-element group 1120: successors 
    -- CP-element group 1120: 	1127 
    -- CP-element group 1120:  members (5) 
      -- CP-element group 1120: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/SplitProtocol/$exit
      -- CP-element group 1120: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/type_cast_3804/$exit
      -- CP-element group 1120: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_sources/$exit
      -- CP-element group 1120: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/$exit
      -- CP-element group 1120: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3801/phi_stmt_3801_req
      -- 
    phi_stmt_3801_req_13080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3801_req_13080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1120), ack => phi_stmt_3801_req_0); -- 
    zeropad3D_cp_element_group_1120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1118) & zeropad3D_CP_2067_elements(1119);
      gj_zeropad3D_cp_element_group_1120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1121:  transition  input  bypass 
    -- CP-element group 1121: predecessors 
    -- CP-element group 1121: 	579 
    -- CP-element group 1121: successors 
    -- CP-element group 1121: 	1123 
    -- CP-element group 1121:  members (2) 
      -- CP-element group 1121: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/Sample/$exit
      -- CP-element group 1121: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/Sample/ra
      -- 
    ra_13097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3811_inst_ack_0, ack => zeropad3D_CP_2067_elements(1121)); -- 
    -- CP-element group 1122:  transition  input  bypass 
    -- CP-element group 1122: predecessors 
    -- CP-element group 1122: 	579 
    -- CP-element group 1122: successors 
    -- CP-element group 1122: 	1123 
    -- CP-element group 1122:  members (2) 
      -- CP-element group 1122: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/Update/$exit
      -- CP-element group 1122: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/Update/ca
      -- 
    ca_13102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3811_inst_ack_1, ack => zeropad3D_CP_2067_elements(1122)); -- 
    -- CP-element group 1123:  join  transition  output  bypass 
    -- CP-element group 1123: predecessors 
    -- CP-element group 1123: 	1121 
    -- CP-element group 1123: 	1122 
    -- CP-element group 1123: successors 
    -- CP-element group 1123: 	1127 
    -- CP-element group 1123:  members (5) 
      -- CP-element group 1123: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/$exit
      -- CP-element group 1123: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/$exit
      -- CP-element group 1123: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/$exit
      -- CP-element group 1123: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_sources/type_cast_3811/SplitProtocol/$exit
      -- CP-element group 1123: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3808/phi_stmt_3808_req
      -- 
    phi_stmt_3808_req_13103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3808_req_13103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1123), ack => phi_stmt_3808_req_0); -- 
    zeropad3D_cp_element_group_1123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1121) & zeropad3D_CP_2067_elements(1122);
      gj_zeropad3D_cp_element_group_1123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1124:  transition  input  bypass 
    -- CP-element group 1124: predecessors 
    -- CP-element group 1124: 	579 
    -- CP-element group 1124: successors 
    -- CP-element group 1124: 	1126 
    -- CP-element group 1124:  members (2) 
      -- CP-element group 1124: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/Sample/$exit
      -- CP-element group 1124: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/Sample/ra
      -- 
    ra_13120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3817_inst_ack_0, ack => zeropad3D_CP_2067_elements(1124)); -- 
    -- CP-element group 1125:  transition  input  bypass 
    -- CP-element group 1125: predecessors 
    -- CP-element group 1125: 	579 
    -- CP-element group 1125: successors 
    -- CP-element group 1125: 	1126 
    -- CP-element group 1125:  members (2) 
      -- CP-element group 1125: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/Update/$exit
      -- CP-element group 1125: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/Update/ca
      -- 
    ca_13125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3817_inst_ack_1, ack => zeropad3D_CP_2067_elements(1125)); -- 
    -- CP-element group 1126:  join  transition  output  bypass 
    -- CP-element group 1126: predecessors 
    -- CP-element group 1126: 	1124 
    -- CP-element group 1126: 	1125 
    -- CP-element group 1126: successors 
    -- CP-element group 1126: 	1127 
    -- CP-element group 1126:  members (5) 
      -- CP-element group 1126: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/$exit
      -- CP-element group 1126: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/$exit
      -- CP-element group 1126: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/$exit
      -- CP-element group 1126: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_sources/type_cast_3817/SplitProtocol/$exit
      -- CP-element group 1126: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/phi_stmt_3814/phi_stmt_3814_req
      -- 
    phi_stmt_3814_req_13126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3814_req_13126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1126), ack => phi_stmt_3814_req_0); -- 
    zeropad3D_cp_element_group_1126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1124) & zeropad3D_CP_2067_elements(1125);
      gj_zeropad3D_cp_element_group_1126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1127:  join  transition  bypass 
    -- CP-element group 1127: predecessors 
    -- CP-element group 1127: 	1120 
    -- CP-element group 1127: 	1123 
    -- CP-element group 1127: 	1126 
    -- CP-element group 1127: successors 
    -- CP-element group 1127: 	1128 
    -- CP-element group 1127:  members (1) 
      -- CP-element group 1127: 	 branch_block_stmt_655/ifx_xthen1227_ifx_xend1269_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1120) & zeropad3D_CP_2067_elements(1123) & zeropad3D_CP_2067_elements(1126);
      gj_zeropad3D_cp_element_group_1127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1128:  merge  fork  transition  place  bypass 
    -- CP-element group 1128: predecessors 
    -- CP-element group 1128: 	1117 
    -- CP-element group 1128: 	1127 
    -- CP-element group 1128: successors 
    -- CP-element group 1128: 	1129 
    -- CP-element group 1128: 	1130 
    -- CP-element group 1128: 	1131 
    -- CP-element group 1128:  members (2) 
      -- CP-element group 1128: 	 branch_block_stmt_655/merge_stmt_3800_PhiReqMerge
      -- CP-element group 1128: 	 branch_block_stmt_655/merge_stmt_3800_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1128) <= OrReduce(zeropad3D_CP_2067_elements(1117) & zeropad3D_CP_2067_elements(1127));
    -- CP-element group 1129:  transition  input  bypass 
    -- CP-element group 1129: predecessors 
    -- CP-element group 1129: 	1128 
    -- CP-element group 1129: successors 
    -- CP-element group 1129: 	1132 
    -- CP-element group 1129:  members (1) 
      -- CP-element group 1129: 	 branch_block_stmt_655/merge_stmt_3800_PhiAck/phi_stmt_3801_ack
      -- 
    phi_stmt_3801_ack_13131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3801_ack_0, ack => zeropad3D_CP_2067_elements(1129)); -- 
    -- CP-element group 1130:  transition  input  bypass 
    -- CP-element group 1130: predecessors 
    -- CP-element group 1130: 	1128 
    -- CP-element group 1130: successors 
    -- CP-element group 1130: 	1132 
    -- CP-element group 1130:  members (1) 
      -- CP-element group 1130: 	 branch_block_stmt_655/merge_stmt_3800_PhiAck/phi_stmt_3808_ack
      -- 
    phi_stmt_3808_ack_13132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3808_ack_0, ack => zeropad3D_CP_2067_elements(1130)); -- 
    -- CP-element group 1131:  transition  input  bypass 
    -- CP-element group 1131: predecessors 
    -- CP-element group 1131: 	1128 
    -- CP-element group 1131: successors 
    -- CP-element group 1131: 	1132 
    -- CP-element group 1131:  members (1) 
      -- CP-element group 1131: 	 branch_block_stmt_655/merge_stmt_3800_PhiAck/phi_stmt_3814_ack
      -- 
    phi_stmt_3814_ack_13133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3814_ack_0, ack => zeropad3D_CP_2067_elements(1131)); -- 
    -- CP-element group 1132:  join  transition  bypass 
    -- CP-element group 1132: predecessors 
    -- CP-element group 1132: 	1129 
    -- CP-element group 1132: 	1130 
    -- CP-element group 1132: 	1131 
    -- CP-element group 1132: successors 
    -- CP-element group 1132: 	6 
    -- CP-element group 1132:  members (1) 
      -- CP-element group 1132: 	 branch_block_stmt_655/merge_stmt_3800_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1132: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1132"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1129) & zeropad3D_CP_2067_elements(1130) & zeropad3D_CP_2067_elements(1131);
      gj_zeropad3D_cp_element_group_1132 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1133:  transition  input  bypass 
    -- CP-element group 1133: predecessors 
    -- CP-element group 1133: 	597 
    -- CP-element group 1133: successors 
    -- CP-element group 1133: 	1135 
    -- CP-element group 1133:  members (2) 
      -- CP-element group 1133: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/Sample/$exit
      -- CP-element group 1133: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/Sample/ra
      -- 
    ra_13153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3826_inst_ack_0, ack => zeropad3D_CP_2067_elements(1133)); -- 
    -- CP-element group 1134:  transition  input  bypass 
    -- CP-element group 1134: predecessors 
    -- CP-element group 1134: 	597 
    -- CP-element group 1134: successors 
    -- CP-element group 1134: 	1135 
    -- CP-element group 1134:  members (2) 
      -- CP-element group 1134: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/Update/$exit
      -- CP-element group 1134: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/Update/ca
      -- 
    ca_13158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3826_inst_ack_1, ack => zeropad3D_CP_2067_elements(1134)); -- 
    -- CP-element group 1135:  join  transition  output  bypass 
    -- CP-element group 1135: predecessors 
    -- CP-element group 1135: 	1133 
    -- CP-element group 1135: 	1134 
    -- CP-element group 1135: successors 
    -- CP-element group 1135: 	1139 
    -- CP-element group 1135:  members (5) 
      -- CP-element group 1135: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/$exit
      -- CP-element group 1135: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/$exit
      -- CP-element group 1135: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/$exit
      -- CP-element group 1135: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_sources/type_cast_3826/SplitProtocol/$exit
      -- CP-element group 1135: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3823/phi_stmt_3823_req
      -- 
    phi_stmt_3823_req_13159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3823_req_13159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1135), ack => phi_stmt_3823_req_0); -- 
    zeropad3D_cp_element_group_1135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1133) & zeropad3D_CP_2067_elements(1134);
      gj_zeropad3D_cp_element_group_1135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1136:  transition  input  bypass 
    -- CP-element group 1136: predecessors 
    -- CP-element group 1136: 	597 
    -- CP-element group 1136: successors 
    -- CP-element group 1136: 	1138 
    -- CP-element group 1136:  members (2) 
      -- CP-element group 1136: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/Sample/$exit
      -- CP-element group 1136: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/Sample/ra
      -- 
    ra_13176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3830_inst_ack_0, ack => zeropad3D_CP_2067_elements(1136)); -- 
    -- CP-element group 1137:  transition  input  bypass 
    -- CP-element group 1137: predecessors 
    -- CP-element group 1137: 	597 
    -- CP-element group 1137: successors 
    -- CP-element group 1137: 	1138 
    -- CP-element group 1137:  members (2) 
      -- CP-element group 1137: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/Update/$exit
      -- CP-element group 1137: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/Update/ca
      -- 
    ca_13181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3830_inst_ack_1, ack => zeropad3D_CP_2067_elements(1137)); -- 
    -- CP-element group 1138:  join  transition  output  bypass 
    -- CP-element group 1138: predecessors 
    -- CP-element group 1138: 	1136 
    -- CP-element group 1138: 	1137 
    -- CP-element group 1138: successors 
    -- CP-element group 1138: 	1139 
    -- CP-element group 1138:  members (5) 
      -- CP-element group 1138: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/$exit
      -- CP-element group 1138: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/$exit
      -- CP-element group 1138: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/$exit
      -- CP-element group 1138: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_sources/type_cast_3830/SplitProtocol/$exit
      -- CP-element group 1138: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/phi_stmt_3827/phi_stmt_3827_req
      -- 
    phi_stmt_3827_req_13182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3827_req_13182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1138), ack => phi_stmt_3827_req_0); -- 
    zeropad3D_cp_element_group_1138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1136) & zeropad3D_CP_2067_elements(1137);
      gj_zeropad3D_cp_element_group_1138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1139:  join  fork  transition  place  bypass 
    -- CP-element group 1139: predecessors 
    -- CP-element group 1139: 	1135 
    -- CP-element group 1139: 	1138 
    -- CP-element group 1139: successors 
    -- CP-element group 1139: 	1140 
    -- CP-element group 1139: 	1141 
    -- CP-element group 1139:  members (3) 
      -- CP-element group 1139: 	 branch_block_stmt_655/ifx_xelse1232_whilex_xend1270_PhiReq/$exit
      -- CP-element group 1139: 	 branch_block_stmt_655/merge_stmt_3822_PhiReqMerge
      -- CP-element group 1139: 	 branch_block_stmt_655/merge_stmt_3822_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_1139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1135) & zeropad3D_CP_2067_elements(1138);
      gj_zeropad3D_cp_element_group_1139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1140:  transition  input  bypass 
    -- CP-element group 1140: predecessors 
    -- CP-element group 1140: 	1139 
    -- CP-element group 1140: successors 
    -- CP-element group 1140: 	1142 
    -- CP-element group 1140:  members (1) 
      -- CP-element group 1140: 	 branch_block_stmt_655/merge_stmt_3822_PhiAck/phi_stmt_3823_ack
      -- 
    phi_stmt_3823_ack_13187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3823_ack_0, ack => zeropad3D_CP_2067_elements(1140)); -- 
    -- CP-element group 1141:  transition  input  bypass 
    -- CP-element group 1141: predecessors 
    -- CP-element group 1141: 	1139 
    -- CP-element group 1141: successors 
    -- CP-element group 1141: 	1142 
    -- CP-element group 1141:  members (1) 
      -- CP-element group 1141: 	 branch_block_stmt_655/merge_stmt_3822_PhiAck/phi_stmt_3827_ack
      -- 
    phi_stmt_3827_ack_13188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3827_ack_0, ack => zeropad3D_CP_2067_elements(1141)); -- 
    -- CP-element group 1142:  join  fork  transition  place  output  bypass 
    -- CP-element group 1142: predecessors 
    -- CP-element group 1142: 	1140 
    -- CP-element group 1142: 	1141 
    -- CP-element group 1142: successors 
    -- CP-element group 1142: 	599 
    -- CP-element group 1142: 	600 
    -- CP-element group 1142: 	601 
    -- CP-element group 1142: 	602 
    -- CP-element group 1142: 	603 
    -- CP-element group 1142: 	604 
    -- CP-element group 1142: 	605 
    -- CP-element group 1142: 	606 
    -- CP-element group 1142: 	607 
    -- CP-element group 1142: 	608 
    -- CP-element group 1142: 	610 
    -- CP-element group 1142: 	612 
    -- CP-element group 1142: 	614 
    -- CP-element group 1142: 	616 
    -- CP-element group 1142: 	618 
    -- CP-element group 1142:  members (73) 
      -- CP-element group 1142: 	 branch_block_stmt_655/merge_stmt_3822__exit__
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925__entry__
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_Update/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_sample_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_Sample/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_Sample/rr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3834_Update/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_sample_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_word_address_calculated
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_root_address_calculated
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Sample/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Sample/word_access_start/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Sample/word_access_start/word_0/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Sample/word_access_start/word_0/rr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/word_access_complete/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/word_access_complete/word_0/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_pad_3849_Update/word_access_complete/word_0/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_sample_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_word_address_calculated
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_root_address_calculated
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Sample/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Sample/word_access_start/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Sample/word_access_start/word_0/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Sample/word_access_start/word_0/rr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/word_access_complete/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/word_access_complete/word_0/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_depth_high_3852_Update/word_access_complete/word_0/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_sample_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_word_address_calculated
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_root_address_calculated
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Sample/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Sample/word_access_start/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Sample/word_access_start/word_0/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Sample/word_access_start/word_0/rr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/word_access_complete/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/word_access_complete/word_0/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_depth_high_3855_Update/word_access_complete/word_0/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_sample_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_word_address_calculated
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_root_address_calculated
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Sample/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Sample/word_access_start/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Sample/word_access_start/word_0/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Sample/word_access_start/word_0/rr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/word_access_complete/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/word_access_complete/word_0/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/LOAD_out_col_high_3858_Update/word_access_complete/word_0/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3862_Update/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3866_Update/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3870_Update/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_Update/$entry
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3879_Update/cr
      -- CP-element group 1142: 	 branch_block_stmt_655/assign_stmt_3835_to_assign_stmt_3925/type_cast_3883_update_start_
      -- CP-element group 1142: 	 branch_block_stmt_655/merge_stmt_3822_PhiAck/$exit
      -- 
    cr_8832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => type_cast_3883_inst_req_1); -- 
    rr_8625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => type_cast_3834_inst_req_0); -- 
    cr_8630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => type_cast_3834_inst_req_1); -- 
    rr_8647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => LOAD_pad_3849_load_0_req_0); -- 
    cr_8658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => LOAD_pad_3849_load_0_req_1); -- 
    rr_8680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => LOAD_depth_high_3852_load_0_req_0); -- 
    cr_8691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => LOAD_depth_high_3852_load_0_req_1); -- 
    rr_8713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => LOAD_out_depth_high_3855_load_0_req_0); -- 
    cr_8724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => LOAD_out_depth_high_3855_load_0_req_1); -- 
    rr_8746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => LOAD_out_col_high_3858_load_0_req_0); -- 
    cr_8757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => LOAD_out_col_high_3858_load_0_req_1); -- 
    cr_8776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => type_cast_3862_inst_req_1); -- 
    cr_8790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => type_cast_3866_inst_req_1); -- 
    cr_8804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => type_cast_3870_inst_req_1); -- 
    cr_8818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1142), ack => type_cast_3879_inst_req_1); -- 
    zeropad3D_cp_element_group_1142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1140) & zeropad3D_CP_2067_elements(1141);
      gj_zeropad3D_cp_element_group_1142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1143:  transition  input  bypass 
    -- CP-element group 1143: predecessors 
    -- CP-element group 1143: 	7 
    -- CP-element group 1143: successors 
    -- CP-element group 1143: 	1145 
    -- CP-element group 1143:  members (2) 
      -- CP-element group 1143: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/Sample/$exit
      -- CP-element group 1143: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/Sample/ra
      -- 
    ra_13208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3934_inst_ack_0, ack => zeropad3D_CP_2067_elements(1143)); -- 
    -- CP-element group 1144:  transition  input  bypass 
    -- CP-element group 1144: predecessors 
    -- CP-element group 1144: 	7 
    -- CP-element group 1144: successors 
    -- CP-element group 1144: 	1145 
    -- CP-element group 1144:  members (2) 
      -- CP-element group 1144: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/Update/$exit
      -- CP-element group 1144: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/Update/ca
      -- 
    ca_13213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3934_inst_ack_1, ack => zeropad3D_CP_2067_elements(1144)); -- 
    -- CP-element group 1145:  join  transition  output  bypass 
    -- CP-element group 1145: predecessors 
    -- CP-element group 1145: 	1143 
    -- CP-element group 1145: 	1144 
    -- CP-element group 1145: successors 
    -- CP-element group 1145: 	1152 
    -- CP-element group 1145:  members (5) 
      -- CP-element group 1145: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/$exit
      -- CP-element group 1145: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/$exit
      -- CP-element group 1145: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/$exit
      -- CP-element group 1145: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3934/SplitProtocol/$exit
      -- CP-element group 1145: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_req
      -- 
    phi_stmt_3928_req_13214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3928_req_13214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1145), ack => phi_stmt_3928_req_1); -- 
    zeropad3D_cp_element_group_1145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1143) & zeropad3D_CP_2067_elements(1144);
      gj_zeropad3D_cp_element_group_1145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1146:  transition  input  bypass 
    -- CP-element group 1146: predecessors 
    -- CP-element group 1146: 	7 
    -- CP-element group 1146: successors 
    -- CP-element group 1146: 	1148 
    -- CP-element group 1146:  members (2) 
      -- CP-element group 1146: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/Sample/$exit
      -- CP-element group 1146: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/Sample/ra
      -- 
    ra_13231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3938_inst_ack_0, ack => zeropad3D_CP_2067_elements(1146)); -- 
    -- CP-element group 1147:  transition  input  bypass 
    -- CP-element group 1147: predecessors 
    -- CP-element group 1147: 	7 
    -- CP-element group 1147: successors 
    -- CP-element group 1147: 	1148 
    -- CP-element group 1147:  members (2) 
      -- CP-element group 1147: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/Update/$exit
      -- CP-element group 1147: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/Update/ca
      -- 
    ca_13236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3938_inst_ack_1, ack => zeropad3D_CP_2067_elements(1147)); -- 
    -- CP-element group 1148:  join  transition  output  bypass 
    -- CP-element group 1148: predecessors 
    -- CP-element group 1148: 	1146 
    -- CP-element group 1148: 	1147 
    -- CP-element group 1148: successors 
    -- CP-element group 1148: 	1152 
    -- CP-element group 1148:  members (5) 
      -- CP-element group 1148: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/$exit
      -- CP-element group 1148: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/$exit
      -- CP-element group 1148: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/$exit
      -- CP-element group 1148: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3938/SplitProtocol/$exit
      -- CP-element group 1148: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_req
      -- 
    phi_stmt_3935_req_13237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3935_req_13237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1148), ack => phi_stmt_3935_req_0); -- 
    zeropad3D_cp_element_group_1148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1146) & zeropad3D_CP_2067_elements(1147);
      gj_zeropad3D_cp_element_group_1148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1149:  transition  input  bypass 
    -- CP-element group 1149: predecessors 
    -- CP-element group 1149: 	7 
    -- CP-element group 1149: successors 
    -- CP-element group 1149: 	1151 
    -- CP-element group 1149:  members (2) 
      -- CP-element group 1149: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/Sample/$exit
      -- CP-element group 1149: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/Sample/ra
      -- 
    ra_13254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3947_inst_ack_0, ack => zeropad3D_CP_2067_elements(1149)); -- 
    -- CP-element group 1150:  transition  input  bypass 
    -- CP-element group 1150: predecessors 
    -- CP-element group 1150: 	7 
    -- CP-element group 1150: successors 
    -- CP-element group 1150: 	1151 
    -- CP-element group 1150:  members (2) 
      -- CP-element group 1150: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/Update/$exit
      -- CP-element group 1150: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/Update/ca
      -- 
    ca_13259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3947_inst_ack_1, ack => zeropad3D_CP_2067_elements(1150)); -- 
    -- CP-element group 1151:  join  transition  output  bypass 
    -- CP-element group 1151: predecessors 
    -- CP-element group 1151: 	1149 
    -- CP-element group 1151: 	1150 
    -- CP-element group 1151: successors 
    -- CP-element group 1151: 	1152 
    -- CP-element group 1151:  members (5) 
      -- CP-element group 1151: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/$exit
      -- CP-element group 1151: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/$exit
      -- CP-element group 1151: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/$exit
      -- CP-element group 1151: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3947/SplitProtocol/$exit
      -- CP-element group 1151: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_req
      -- 
    phi_stmt_3941_req_13260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3941_req_13260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1151), ack => phi_stmt_3941_req_1); -- 
    zeropad3D_cp_element_group_1151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1149) & zeropad3D_CP_2067_elements(1150);
      gj_zeropad3D_cp_element_group_1151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1152:  join  transition  bypass 
    -- CP-element group 1152: predecessors 
    -- CP-element group 1152: 	1145 
    -- CP-element group 1152: 	1148 
    -- CP-element group 1152: 	1151 
    -- CP-element group 1152: successors 
    -- CP-element group 1152: 	1159 
    -- CP-element group 1152:  members (1) 
      -- CP-element group 1152: 	 branch_block_stmt_655/ifx_xend1486_whilex_xbody1331_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1152: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1152"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1145) & zeropad3D_CP_2067_elements(1148) & zeropad3D_CP_2067_elements(1151);
      gj_zeropad3D_cp_element_group_1152 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1153:  transition  output  delay-element  bypass 
    -- CP-element group 1153: predecessors 
    -- CP-element group 1153: 	619 
    -- CP-element group 1153: successors 
    -- CP-element group 1153: 	1158 
    -- CP-element group 1153:  members (4) 
      -- CP-element group 1153: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3928/$exit
      -- CP-element group 1153: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/$exit
      -- CP-element group 1153: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_sources/type_cast_3932_konst_delay_trans
      -- CP-element group 1153: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3928/phi_stmt_3928_req
      -- 
    phi_stmt_3928_req_13271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3928_req_13271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1153), ack => phi_stmt_3928_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(1153) is a control-delay.
    cp_element_1153_delay: control_delay_element  generic map(name => " 1153_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(619), ack => zeropad3D_CP_2067_elements(1153), clk => clk, reset =>reset);
    -- CP-element group 1154:  transition  input  bypass 
    -- CP-element group 1154: predecessors 
    -- CP-element group 1154: 	619 
    -- CP-element group 1154: successors 
    -- CP-element group 1154: 	1156 
    -- CP-element group 1154:  members (2) 
      -- CP-element group 1154: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/Sample/$exit
      -- CP-element group 1154: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/Sample/ra
      -- 
    ra_13288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3940_inst_ack_0, ack => zeropad3D_CP_2067_elements(1154)); -- 
    -- CP-element group 1155:  transition  input  bypass 
    -- CP-element group 1155: predecessors 
    -- CP-element group 1155: 	619 
    -- CP-element group 1155: successors 
    -- CP-element group 1155: 	1156 
    -- CP-element group 1155:  members (2) 
      -- CP-element group 1155: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/Update/$exit
      -- CP-element group 1155: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/Update/ca
      -- 
    ca_13293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3940_inst_ack_1, ack => zeropad3D_CP_2067_elements(1155)); -- 
    -- CP-element group 1156:  join  transition  output  bypass 
    -- CP-element group 1156: predecessors 
    -- CP-element group 1156: 	1154 
    -- CP-element group 1156: 	1155 
    -- CP-element group 1156: successors 
    -- CP-element group 1156: 	1158 
    -- CP-element group 1156:  members (5) 
      -- CP-element group 1156: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/$exit
      -- CP-element group 1156: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/$exit
      -- CP-element group 1156: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/$exit
      -- CP-element group 1156: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_sources/type_cast_3940/SplitProtocol/$exit
      -- CP-element group 1156: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3935/phi_stmt_3935_req
      -- 
    phi_stmt_3935_req_13294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3935_req_13294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1156), ack => phi_stmt_3935_req_1); -- 
    zeropad3D_cp_element_group_1156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1154) & zeropad3D_CP_2067_elements(1155);
      gj_zeropad3D_cp_element_group_1156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1157:  transition  output  delay-element  bypass 
    -- CP-element group 1157: predecessors 
    -- CP-element group 1157: 	619 
    -- CP-element group 1157: successors 
    -- CP-element group 1157: 	1158 
    -- CP-element group 1157:  members (4) 
      -- CP-element group 1157: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3941/$exit
      -- CP-element group 1157: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/$exit
      -- CP-element group 1157: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_sources/type_cast_3945_konst_delay_trans
      -- CP-element group 1157: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/phi_stmt_3941/phi_stmt_3941_req
      -- 
    phi_stmt_3941_req_13302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3941_req_13302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1157), ack => phi_stmt_3941_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(1157) is a control-delay.
    cp_element_1157_delay: control_delay_element  generic map(name => " 1157_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(619), ack => zeropad3D_CP_2067_elements(1157), clk => clk, reset =>reset);
    -- CP-element group 1158:  join  transition  bypass 
    -- CP-element group 1158: predecessors 
    -- CP-element group 1158: 	1153 
    -- CP-element group 1158: 	1156 
    -- CP-element group 1158: 	1157 
    -- CP-element group 1158: successors 
    -- CP-element group 1158: 	1159 
    -- CP-element group 1158:  members (1) 
      -- CP-element group 1158: 	 branch_block_stmt_655/whilex_xend1270_whilex_xbody1331_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1153) & zeropad3D_CP_2067_elements(1156) & zeropad3D_CP_2067_elements(1157);
      gj_zeropad3D_cp_element_group_1158 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1159:  merge  fork  transition  place  bypass 
    -- CP-element group 1159: predecessors 
    -- CP-element group 1159: 	1152 
    -- CP-element group 1159: 	1158 
    -- CP-element group 1159: successors 
    -- CP-element group 1159: 	1160 
    -- CP-element group 1159: 	1161 
    -- CP-element group 1159: 	1162 
    -- CP-element group 1159:  members (2) 
      -- CP-element group 1159: 	 branch_block_stmt_655/merge_stmt_3927_PhiReqMerge
      -- CP-element group 1159: 	 branch_block_stmt_655/merge_stmt_3927_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1159) <= OrReduce(zeropad3D_CP_2067_elements(1152) & zeropad3D_CP_2067_elements(1158));
    -- CP-element group 1160:  transition  input  bypass 
    -- CP-element group 1160: predecessors 
    -- CP-element group 1160: 	1159 
    -- CP-element group 1160: successors 
    -- CP-element group 1160: 	1163 
    -- CP-element group 1160:  members (1) 
      -- CP-element group 1160: 	 branch_block_stmt_655/merge_stmt_3927_PhiAck/phi_stmt_3928_ack
      -- 
    phi_stmt_3928_ack_13307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3928_ack_0, ack => zeropad3D_CP_2067_elements(1160)); -- 
    -- CP-element group 1161:  transition  input  bypass 
    -- CP-element group 1161: predecessors 
    -- CP-element group 1161: 	1159 
    -- CP-element group 1161: successors 
    -- CP-element group 1161: 	1163 
    -- CP-element group 1161:  members (1) 
      -- CP-element group 1161: 	 branch_block_stmt_655/merge_stmt_3927_PhiAck/phi_stmt_3935_ack
      -- 
    phi_stmt_3935_ack_13308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3935_ack_0, ack => zeropad3D_CP_2067_elements(1161)); -- 
    -- CP-element group 1162:  transition  input  bypass 
    -- CP-element group 1162: predecessors 
    -- CP-element group 1162: 	1159 
    -- CP-element group 1162: successors 
    -- CP-element group 1162: 	1163 
    -- CP-element group 1162:  members (1) 
      -- CP-element group 1162: 	 branch_block_stmt_655/merge_stmt_3927_PhiAck/phi_stmt_3941_ack
      -- 
    phi_stmt_3941_ack_13309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3941_ack_0, ack => zeropad3D_CP_2067_elements(1162)); -- 
    -- CP-element group 1163:  join  fork  transition  place  output  bypass 
    -- CP-element group 1163: predecessors 
    -- CP-element group 1163: 	1160 
    -- CP-element group 1163: 	1161 
    -- CP-element group 1163: 	1162 
    -- CP-element group 1163: successors 
    -- CP-element group 1163: 	620 
    -- CP-element group 1163: 	621 
    -- CP-element group 1163:  members (10) 
      -- CP-element group 1163: 	 branch_block_stmt_655/merge_stmt_3927__exit__
      -- CP-element group 1163: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960__entry__
      -- CP-element group 1163: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/$entry
      -- CP-element group 1163: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_sample_start_
      -- CP-element group 1163: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_Update/cr
      -- CP-element group 1163: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_Update/$entry
      -- CP-element group 1163: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_Sample/rr
      -- CP-element group 1163: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_Sample/$entry
      -- CP-element group 1163: 	 branch_block_stmt_655/assign_stmt_3953_to_assign_stmt_3960/type_cast_3952_update_start_
      -- CP-element group 1163: 	 branch_block_stmt_655/merge_stmt_3927_PhiAck/$exit
      -- 
    cr_8849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1163), ack => type_cast_3952_inst_req_1); -- 
    rr_8844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1163), ack => type_cast_3952_inst_req_0); -- 
    zeropad3D_cp_element_group_1163: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1163"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1160) & zeropad3D_CP_2067_elements(1161) & zeropad3D_CP_2067_elements(1162);
      gj_zeropad3D_cp_element_group_1163 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1164:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1164: predecessors 
    -- CP-element group 1164: 	622 
    -- CP-element group 1164: 	629 
    -- CP-element group 1164: 	632 
    -- CP-element group 1164: 	639 
    -- CP-element group 1164: successors 
    -- CP-element group 1164: 	640 
    -- CP-element group 1164: 	641 
    -- CP-element group 1164: 	642 
    -- CP-element group 1164: 	643 
    -- CP-element group 1164: 	646 
    -- CP-element group 1164: 	648 
    -- CP-element group 1164: 	650 
    -- CP-element group 1164: 	652 
    -- CP-element group 1164:  members (33) 
      -- CP-element group 1164: 	 branch_block_stmt_655/merge_stmt_4044__exit__
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100__entry__
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_Update/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_Update/cr
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_Sample/rr
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_Sample/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_update_start_
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_complete/req
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/addr_of_4094_complete/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_update_start_
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_Update/cr
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_Update/req
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_Update/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4048_sample_start_
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Update/word_access_complete/word_0/cr
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Update/word_access_complete/word_0/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_Update/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4087_update_start_
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Update/word_access_complete/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_Update/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_Update/cr
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/array_obj_ref_4093_final_index_sum_regn_update_start
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_Update/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_Sample/rr
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_Sample/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_update_start_
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/type_cast_4053_sample_start_
      -- CP-element group 1164: 	 branch_block_stmt_655/assign_stmt_4049_to_assign_stmt_4100/ptr_deref_4097_update_start_
      -- CP-element group 1164: 	 branch_block_stmt_655/merge_stmt_4044_PhiReqMerge
      -- CP-element group 1164: 	 branch_block_stmt_655/merge_stmt_4044_PhiAck/$entry
      -- CP-element group 1164: 	 branch_block_stmt_655/merge_stmt_4044_PhiAck/$exit
      -- CP-element group 1164: 	 branch_block_stmt_655/merge_stmt_4044_PhiAck/dummy
      -- 
    cr_9059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1164), ack => type_cast_4048_inst_req_1); -- 
    rr_9054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1164), ack => type_cast_4048_inst_req_0); -- 
    req_9133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1164), ack => addr_of_4094_final_reg_req_1); -- 
    cr_9087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1164), ack => type_cast_4087_inst_req_1); -- 
    req_9118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1164), ack => array_obj_ref_4093_index_offset_req_1); -- 
    cr_9183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1164), ack => ptr_deref_4097_store_0_req_1); -- 
    cr_9073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1164), ack => type_cast_4053_inst_req_1); -- 
    rr_9068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1164), ack => type_cast_4053_inst_req_0); -- 
    zeropad3D_CP_2067_elements(1164) <= OrReduce(zeropad3D_CP_2067_elements(622) & zeropad3D_CP_2067_elements(629) & zeropad3D_CP_2067_elements(632) & zeropad3D_CP_2067_elements(639));
    -- CP-element group 1165:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1165: predecessors 
    -- CP-element group 1165: 	653 
    -- CP-element group 1165: 	673 
    -- CP-element group 1165: successors 
    -- CP-element group 1165: 	674 
    -- CP-element group 1165: 	675 
    -- CP-element group 1165:  members (13) 
      -- CP-element group 1165: 	 branch_block_stmt_655/merge_stmt_4209__exit__
      -- CP-element group 1165: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227__entry__
      -- CP-element group 1165: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/$entry
      -- CP-element group 1165: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_sample_start_
      -- CP-element group 1165: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_update_start_
      -- CP-element group 1165: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_Sample/$entry
      -- CP-element group 1165: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_Sample/rr
      -- CP-element group 1165: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_Update/$entry
      -- CP-element group 1165: 	 branch_block_stmt_655/assign_stmt_4214_to_assign_stmt_4227/type_cast_4213_Update/cr
      -- CP-element group 1165: 	 branch_block_stmt_655/merge_stmt_4209_PhiReqMerge
      -- CP-element group 1165: 	 branch_block_stmt_655/merge_stmt_4209_PhiAck/$entry
      -- CP-element group 1165: 	 branch_block_stmt_655/merge_stmt_4209_PhiAck/$exit
      -- CP-element group 1165: 	 branch_block_stmt_655/merge_stmt_4209_PhiAck/dummy
      -- 
    rr_9432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1165), ack => type_cast_4213_inst_req_0); -- 
    cr_9437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1165), ack => type_cast_4213_inst_req_1); -- 
    zeropad3D_CP_2067_elements(1165) <= OrReduce(zeropad3D_CP_2067_elements(653) & zeropad3D_CP_2067_elements(673));
    -- CP-element group 1166:  transition  output  delay-element  bypass 
    -- CP-element group 1166: predecessors 
    -- CP-element group 1166: 	695 
    -- CP-element group 1166: successors 
    -- CP-element group 1166: 	1173 
    -- CP-element group 1166:  members (4) 
      -- CP-element group 1166: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4322/$exit
      -- CP-element group 1166: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/$exit
      -- CP-element group 1166: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4328_konst_delay_trans
      -- CP-element group 1166: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_req
      -- 
    phi_stmt_4322_req_13420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4322_req_13420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1166), ack => phi_stmt_4322_req_1); -- 
    -- Element group zeropad3D_CP_2067_elements(1166) is a control-delay.
    cp_element_1166_delay: control_delay_element  generic map(name => " 1166_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(695), ack => zeropad3D_CP_2067_elements(1166), clk => clk, reset =>reset);
    -- CP-element group 1167:  transition  input  bypass 
    -- CP-element group 1167: predecessors 
    -- CP-element group 1167: 	695 
    -- CP-element group 1167: successors 
    -- CP-element group 1167: 	1169 
    -- CP-element group 1167:  members (2) 
      -- CP-element group 1167: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/Sample/$exit
      -- CP-element group 1167: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/Sample/ra
      -- 
    ra_13437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4334_inst_ack_0, ack => zeropad3D_CP_2067_elements(1167)); -- 
    -- CP-element group 1168:  transition  input  bypass 
    -- CP-element group 1168: predecessors 
    -- CP-element group 1168: 	695 
    -- CP-element group 1168: successors 
    -- CP-element group 1168: 	1169 
    -- CP-element group 1168:  members (2) 
      -- CP-element group 1168: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/Update/$exit
      -- CP-element group 1168: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/Update/ca
      -- 
    ca_13442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4334_inst_ack_1, ack => zeropad3D_CP_2067_elements(1168)); -- 
    -- CP-element group 1169:  join  transition  output  bypass 
    -- CP-element group 1169: predecessors 
    -- CP-element group 1169: 	1167 
    -- CP-element group 1169: 	1168 
    -- CP-element group 1169: successors 
    -- CP-element group 1169: 	1173 
    -- CP-element group 1169:  members (5) 
      -- CP-element group 1169: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/$exit
      -- CP-element group 1169: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/$exit
      -- CP-element group 1169: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/$exit
      -- CP-element group 1169: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4334/SplitProtocol/$exit
      -- CP-element group 1169: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_req
      -- 
    phi_stmt_4329_req_13443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4329_req_13443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1169), ack => phi_stmt_4329_req_1); -- 
    zeropad3D_cp_element_group_1169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1167) & zeropad3D_CP_2067_elements(1168);
      gj_zeropad3D_cp_element_group_1169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1170:  transition  input  bypass 
    -- CP-element group 1170: predecessors 
    -- CP-element group 1170: 	695 
    -- CP-element group 1170: successors 
    -- CP-element group 1170: 	1172 
    -- CP-element group 1170:  members (2) 
      -- CP-element group 1170: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/Sample/$exit
      -- CP-element group 1170: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/Sample/ra
      -- 
    ra_13460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4340_inst_ack_0, ack => zeropad3D_CP_2067_elements(1170)); -- 
    -- CP-element group 1171:  transition  input  bypass 
    -- CP-element group 1171: predecessors 
    -- CP-element group 1171: 	695 
    -- CP-element group 1171: successors 
    -- CP-element group 1171: 	1172 
    -- CP-element group 1171:  members (2) 
      -- CP-element group 1171: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/Update/$exit
      -- CP-element group 1171: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/Update/ca
      -- 
    ca_13465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4340_inst_ack_1, ack => zeropad3D_CP_2067_elements(1171)); -- 
    -- CP-element group 1172:  join  transition  output  bypass 
    -- CP-element group 1172: predecessors 
    -- CP-element group 1172: 	1170 
    -- CP-element group 1172: 	1171 
    -- CP-element group 1172: successors 
    -- CP-element group 1172: 	1173 
    -- CP-element group 1172:  members (5) 
      -- CP-element group 1172: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/$exit
      -- CP-element group 1172: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/$exit
      -- CP-element group 1172: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/$exit
      -- CP-element group 1172: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4340/SplitProtocol/$exit
      -- CP-element group 1172: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_req
      -- 
    phi_stmt_4335_req_13466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4335_req_13466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1172), ack => phi_stmt_4335_req_1); -- 
    zeropad3D_cp_element_group_1172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1170) & zeropad3D_CP_2067_elements(1171);
      gj_zeropad3D_cp_element_group_1172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1173:  join  transition  bypass 
    -- CP-element group 1173: predecessors 
    -- CP-element group 1173: 	1166 
    -- CP-element group 1173: 	1169 
    -- CP-element group 1173: 	1172 
    -- CP-element group 1173: successors 
    -- CP-element group 1173: 	1184 
    -- CP-element group 1173:  members (1) 
      -- CP-element group 1173: 	 branch_block_stmt_655/ifx_xelse1450_ifx_xend1486_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1166) & zeropad3D_CP_2067_elements(1169) & zeropad3D_CP_2067_elements(1172);
      gj_zeropad3D_cp_element_group_1173 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1174:  transition  input  bypass 
    -- CP-element group 1174: predecessors 
    -- CP-element group 1174: 	676 
    -- CP-element group 1174: successors 
    -- CP-element group 1174: 	1176 
    -- CP-element group 1174:  members (2) 
      -- CP-element group 1174: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/Sample/$exit
      -- CP-element group 1174: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/Sample/ra
      -- 
    ra_13486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4325_inst_ack_0, ack => zeropad3D_CP_2067_elements(1174)); -- 
    -- CP-element group 1175:  transition  input  bypass 
    -- CP-element group 1175: predecessors 
    -- CP-element group 1175: 	676 
    -- CP-element group 1175: successors 
    -- CP-element group 1175: 	1176 
    -- CP-element group 1175:  members (2) 
      -- CP-element group 1175: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/Update/$exit
      -- CP-element group 1175: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/Update/ca
      -- 
    ca_13491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4325_inst_ack_1, ack => zeropad3D_CP_2067_elements(1175)); -- 
    -- CP-element group 1176:  join  transition  output  bypass 
    -- CP-element group 1176: predecessors 
    -- CP-element group 1176: 	1174 
    -- CP-element group 1176: 	1175 
    -- CP-element group 1176: successors 
    -- CP-element group 1176: 	1183 
    -- CP-element group 1176:  members (5) 
      -- CP-element group 1176: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/$exit
      -- CP-element group 1176: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/$exit
      -- CP-element group 1176: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/$exit
      -- CP-element group 1176: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_sources/type_cast_4325/SplitProtocol/$exit
      -- CP-element group 1176: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4322/phi_stmt_4322_req
      -- 
    phi_stmt_4322_req_13492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4322_req_13492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1176), ack => phi_stmt_4322_req_0); -- 
    zeropad3D_cp_element_group_1176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1174) & zeropad3D_CP_2067_elements(1175);
      gj_zeropad3D_cp_element_group_1176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1177:  transition  input  bypass 
    -- CP-element group 1177: predecessors 
    -- CP-element group 1177: 	676 
    -- CP-element group 1177: successors 
    -- CP-element group 1177: 	1179 
    -- CP-element group 1177:  members (2) 
      -- CP-element group 1177: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/Sample/$exit
      -- CP-element group 1177: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/Sample/ra
      -- 
    ra_13509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4332_inst_ack_0, ack => zeropad3D_CP_2067_elements(1177)); -- 
    -- CP-element group 1178:  transition  input  bypass 
    -- CP-element group 1178: predecessors 
    -- CP-element group 1178: 	676 
    -- CP-element group 1178: successors 
    -- CP-element group 1178: 	1179 
    -- CP-element group 1178:  members (2) 
      -- CP-element group 1178: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/Update/$exit
      -- CP-element group 1178: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/Update/ca
      -- 
    ca_13514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4332_inst_ack_1, ack => zeropad3D_CP_2067_elements(1178)); -- 
    -- CP-element group 1179:  join  transition  output  bypass 
    -- CP-element group 1179: predecessors 
    -- CP-element group 1179: 	1177 
    -- CP-element group 1179: 	1178 
    -- CP-element group 1179: successors 
    -- CP-element group 1179: 	1183 
    -- CP-element group 1179:  members (5) 
      -- CP-element group 1179: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/$exit
      -- CP-element group 1179: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/$exit
      -- CP-element group 1179: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/$exit
      -- CP-element group 1179: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_sources/type_cast_4332/SplitProtocol/$exit
      -- CP-element group 1179: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4329/phi_stmt_4329_req
      -- 
    phi_stmt_4329_req_13515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4329_req_13515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1179), ack => phi_stmt_4329_req_0); -- 
    zeropad3D_cp_element_group_1179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1177) & zeropad3D_CP_2067_elements(1178);
      gj_zeropad3D_cp_element_group_1179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1180:  transition  input  bypass 
    -- CP-element group 1180: predecessors 
    -- CP-element group 1180: 	676 
    -- CP-element group 1180: successors 
    -- CP-element group 1180: 	1182 
    -- CP-element group 1180:  members (2) 
      -- CP-element group 1180: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/Sample/$exit
      -- CP-element group 1180: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/Sample/ra
      -- 
    ra_13532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4338_inst_ack_0, ack => zeropad3D_CP_2067_elements(1180)); -- 
    -- CP-element group 1181:  transition  input  bypass 
    -- CP-element group 1181: predecessors 
    -- CP-element group 1181: 	676 
    -- CP-element group 1181: successors 
    -- CP-element group 1181: 	1182 
    -- CP-element group 1181:  members (2) 
      -- CP-element group 1181: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/Update/$exit
      -- CP-element group 1181: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/Update/ca
      -- 
    ca_13537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4338_inst_ack_1, ack => zeropad3D_CP_2067_elements(1181)); -- 
    -- CP-element group 1182:  join  transition  output  bypass 
    -- CP-element group 1182: predecessors 
    -- CP-element group 1182: 	1180 
    -- CP-element group 1182: 	1181 
    -- CP-element group 1182: successors 
    -- CP-element group 1182: 	1183 
    -- CP-element group 1182:  members (5) 
      -- CP-element group 1182: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/$exit
      -- CP-element group 1182: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/$exit
      -- CP-element group 1182: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/$exit
      -- CP-element group 1182: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_sources/type_cast_4338/SplitProtocol/$exit
      -- CP-element group 1182: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/phi_stmt_4335/phi_stmt_4335_req
      -- 
    phi_stmt_4335_req_13538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4335_req_13538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1182), ack => phi_stmt_4335_req_0); -- 
    zeropad3D_cp_element_group_1182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1180) & zeropad3D_CP_2067_elements(1181);
      gj_zeropad3D_cp_element_group_1182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1183:  join  transition  bypass 
    -- CP-element group 1183: predecessors 
    -- CP-element group 1183: 	1176 
    -- CP-element group 1183: 	1179 
    -- CP-element group 1183: 	1182 
    -- CP-element group 1183: successors 
    -- CP-element group 1183: 	1184 
    -- CP-element group 1183:  members (1) 
      -- CP-element group 1183: 	 branch_block_stmt_655/ifx_xthen1445_ifx_xend1486_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1183: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1183"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1176) & zeropad3D_CP_2067_elements(1179) & zeropad3D_CP_2067_elements(1182);
      gj_zeropad3D_cp_element_group_1183 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1184:  merge  fork  transition  place  bypass 
    -- CP-element group 1184: predecessors 
    -- CP-element group 1184: 	1173 
    -- CP-element group 1184: 	1183 
    -- CP-element group 1184: successors 
    -- CP-element group 1184: 	1185 
    -- CP-element group 1184: 	1186 
    -- CP-element group 1184: 	1187 
    -- CP-element group 1184:  members (2) 
      -- CP-element group 1184: 	 branch_block_stmt_655/merge_stmt_4321_PhiReqMerge
      -- CP-element group 1184: 	 branch_block_stmt_655/merge_stmt_4321_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1184) <= OrReduce(zeropad3D_CP_2067_elements(1173) & zeropad3D_CP_2067_elements(1183));
    -- CP-element group 1185:  transition  input  bypass 
    -- CP-element group 1185: predecessors 
    -- CP-element group 1185: 	1184 
    -- CP-element group 1185: successors 
    -- CP-element group 1185: 	1188 
    -- CP-element group 1185:  members (1) 
      -- CP-element group 1185: 	 branch_block_stmt_655/merge_stmt_4321_PhiAck/phi_stmt_4322_ack
      -- 
    phi_stmt_4322_ack_13543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4322_ack_0, ack => zeropad3D_CP_2067_elements(1185)); -- 
    -- CP-element group 1186:  transition  input  bypass 
    -- CP-element group 1186: predecessors 
    -- CP-element group 1186: 	1184 
    -- CP-element group 1186: successors 
    -- CP-element group 1186: 	1188 
    -- CP-element group 1186:  members (1) 
      -- CP-element group 1186: 	 branch_block_stmt_655/merge_stmt_4321_PhiAck/phi_stmt_4329_ack
      -- 
    phi_stmt_4329_ack_13544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4329_ack_0, ack => zeropad3D_CP_2067_elements(1186)); -- 
    -- CP-element group 1187:  transition  input  bypass 
    -- CP-element group 1187: predecessors 
    -- CP-element group 1187: 	1184 
    -- CP-element group 1187: successors 
    -- CP-element group 1187: 	1188 
    -- CP-element group 1187:  members (1) 
      -- CP-element group 1187: 	 branch_block_stmt_655/merge_stmt_4321_PhiAck/phi_stmt_4335_ack
      -- 
    phi_stmt_4335_ack_13545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4335_ack_0, ack => zeropad3D_CP_2067_elements(1187)); -- 
    -- CP-element group 1188:  join  transition  bypass 
    -- CP-element group 1188: predecessors 
    -- CP-element group 1188: 	1185 
    -- CP-element group 1188: 	1186 
    -- CP-element group 1188: 	1187 
    -- CP-element group 1188: successors 
    -- CP-element group 1188: 	7 
    -- CP-element group 1188:  members (1) 
      -- CP-element group 1188: 	 branch_block_stmt_655/merge_stmt_4321_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1188: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1188"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1185) & zeropad3D_CP_2067_elements(1186) & zeropad3D_CP_2067_elements(1187);
      gj_zeropad3D_cp_element_group_1188 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1189:  transition  input  bypass 
    -- CP-element group 1189: predecessors 
    -- CP-element group 1189: 	694 
    -- CP-element group 1189: successors 
    -- CP-element group 1189: 	1191 
    -- CP-element group 1189:  members (2) 
      -- CP-element group 1189: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/Sample/$exit
      -- CP-element group 1189: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/Sample/ra
      -- 
    ra_13565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4347_inst_ack_0, ack => zeropad3D_CP_2067_elements(1189)); -- 
    -- CP-element group 1190:  transition  input  bypass 
    -- CP-element group 1190: predecessors 
    -- CP-element group 1190: 	694 
    -- CP-element group 1190: successors 
    -- CP-element group 1190: 	1191 
    -- CP-element group 1190:  members (2) 
      -- CP-element group 1190: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/Update/$exit
      -- CP-element group 1190: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/Update/ca
      -- 
    ca_13570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4347_inst_ack_1, ack => zeropad3D_CP_2067_elements(1190)); -- 
    -- CP-element group 1191:  join  transition  output  bypass 
    -- CP-element group 1191: predecessors 
    -- CP-element group 1191: 	1189 
    -- CP-element group 1191: 	1190 
    -- CP-element group 1191: successors 
    -- CP-element group 1191: 	1198 
    -- CP-element group 1191:  members (5) 
      -- CP-element group 1191: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/$exit
      -- CP-element group 1191: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/$exit
      -- CP-element group 1191: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/$exit
      -- CP-element group 1191: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_sources/type_cast_4347/SplitProtocol/$exit
      -- CP-element group 1191: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4344/phi_stmt_4344_req
      -- 
    phi_stmt_4344_req_13571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4344_req_13571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1191), ack => phi_stmt_4344_req_0); -- 
    zeropad3D_cp_element_group_1191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1189) & zeropad3D_CP_2067_elements(1190);
      gj_zeropad3D_cp_element_group_1191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1192:  transition  input  bypass 
    -- CP-element group 1192: predecessors 
    -- CP-element group 1192: 	694 
    -- CP-element group 1192: successors 
    -- CP-element group 1192: 	1194 
    -- CP-element group 1192:  members (2) 
      -- CP-element group 1192: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/Sample/$exit
      -- CP-element group 1192: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/Sample/ra
      -- 
    ra_13588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4351_inst_ack_0, ack => zeropad3D_CP_2067_elements(1192)); -- 
    -- CP-element group 1193:  transition  input  bypass 
    -- CP-element group 1193: predecessors 
    -- CP-element group 1193: 	694 
    -- CP-element group 1193: successors 
    -- CP-element group 1193: 	1194 
    -- CP-element group 1193:  members (2) 
      -- CP-element group 1193: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/Update/$exit
      -- CP-element group 1193: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/Update/ca
      -- 
    ca_13593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4351_inst_ack_1, ack => zeropad3D_CP_2067_elements(1193)); -- 
    -- CP-element group 1194:  join  transition  output  bypass 
    -- CP-element group 1194: predecessors 
    -- CP-element group 1194: 	1192 
    -- CP-element group 1194: 	1193 
    -- CP-element group 1194: successors 
    -- CP-element group 1194: 	1198 
    -- CP-element group 1194:  members (5) 
      -- CP-element group 1194: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/$exit
      -- CP-element group 1194: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/$exit
      -- CP-element group 1194: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/$exit
      -- CP-element group 1194: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_sources/type_cast_4351/SplitProtocol/$exit
      -- CP-element group 1194: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4348/phi_stmt_4348_req
      -- 
    phi_stmt_4348_req_13594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4348_req_13594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1194), ack => phi_stmt_4348_req_0); -- 
    zeropad3D_cp_element_group_1194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1192) & zeropad3D_CP_2067_elements(1193);
      gj_zeropad3D_cp_element_group_1194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1195:  transition  input  bypass 
    -- CP-element group 1195: predecessors 
    -- CP-element group 1195: 	694 
    -- CP-element group 1195: successors 
    -- CP-element group 1195: 	1197 
    -- CP-element group 1195:  members (2) 
      -- CP-element group 1195: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Sample/$exit
      -- CP-element group 1195: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Sample/ra
      -- 
    ra_13611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4355_inst_ack_0, ack => zeropad3D_CP_2067_elements(1195)); -- 
    -- CP-element group 1196:  transition  input  bypass 
    -- CP-element group 1196: predecessors 
    -- CP-element group 1196: 	694 
    -- CP-element group 1196: successors 
    -- CP-element group 1196: 	1197 
    -- CP-element group 1196:  members (2) 
      -- CP-element group 1196: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Update/$exit
      -- CP-element group 1196: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/Update/ca
      -- 
    ca_13616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4355_inst_ack_1, ack => zeropad3D_CP_2067_elements(1196)); -- 
    -- CP-element group 1197:  join  transition  output  bypass 
    -- CP-element group 1197: predecessors 
    -- CP-element group 1197: 	1195 
    -- CP-element group 1197: 	1196 
    -- CP-element group 1197: successors 
    -- CP-element group 1197: 	1198 
    -- CP-element group 1197:  members (5) 
      -- CP-element group 1197: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/$exit
      -- CP-element group 1197: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/$exit
      -- CP-element group 1197: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/$exit
      -- CP-element group 1197: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_sources/type_cast_4355/SplitProtocol/$exit
      -- CP-element group 1197: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/phi_stmt_4352/phi_stmt_4352_req
      -- 
    phi_stmt_4352_req_13617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4352_req_13617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1197), ack => phi_stmt_4352_req_0); -- 
    zeropad3D_cp_element_group_1197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1195) & zeropad3D_CP_2067_elements(1196);
      gj_zeropad3D_cp_element_group_1197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1198:  join  fork  transition  place  bypass 
    -- CP-element group 1198: predecessors 
    -- CP-element group 1198: 	1191 
    -- CP-element group 1198: 	1194 
    -- CP-element group 1198: 	1197 
    -- CP-element group 1198: successors 
    -- CP-element group 1198: 	1199 
    -- CP-element group 1198: 	1200 
    -- CP-element group 1198: 	1201 
    -- CP-element group 1198:  members (3) 
      -- CP-element group 1198: 	 branch_block_stmt_655/ifx_xelse1450_whilex_xend1487_PhiReq/$exit
      -- CP-element group 1198: 	 branch_block_stmt_655/merge_stmt_4343_PhiReqMerge
      -- CP-element group 1198: 	 branch_block_stmt_655/merge_stmt_4343_PhiAck/$entry
      -- 
    zeropad3D_cp_element_group_1198: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1198"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1191) & zeropad3D_CP_2067_elements(1194) & zeropad3D_CP_2067_elements(1197);
      gj_zeropad3D_cp_element_group_1198 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1199:  transition  input  bypass 
    -- CP-element group 1199: predecessors 
    -- CP-element group 1199: 	1198 
    -- CP-element group 1199: successors 
    -- CP-element group 1199: 	1202 
    -- CP-element group 1199:  members (1) 
      -- CP-element group 1199: 	 branch_block_stmt_655/merge_stmt_4343_PhiAck/phi_stmt_4344_ack
      -- 
    phi_stmt_4344_ack_13622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4344_ack_0, ack => zeropad3D_CP_2067_elements(1199)); -- 
    -- CP-element group 1200:  transition  input  bypass 
    -- CP-element group 1200: predecessors 
    -- CP-element group 1200: 	1198 
    -- CP-element group 1200: successors 
    -- CP-element group 1200: 	1202 
    -- CP-element group 1200:  members (1) 
      -- CP-element group 1200: 	 branch_block_stmt_655/merge_stmt_4343_PhiAck/phi_stmt_4348_ack
      -- 
    phi_stmt_4348_ack_13623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4348_ack_0, ack => zeropad3D_CP_2067_elements(1200)); -- 
    -- CP-element group 1201:  transition  input  bypass 
    -- CP-element group 1201: predecessors 
    -- CP-element group 1201: 	1198 
    -- CP-element group 1201: successors 
    -- CP-element group 1201: 	1202 
    -- CP-element group 1201:  members (1) 
      -- CP-element group 1201: 	 branch_block_stmt_655/merge_stmt_4343_PhiAck/phi_stmt_4352_ack
      -- 
    phi_stmt_4352_ack_13624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4352_ack_0, ack => zeropad3D_CP_2067_elements(1201)); -- 
    -- CP-element group 1202:  join  fork  transition  place  output  bypass 
    -- CP-element group 1202: predecessors 
    -- CP-element group 1202: 	1199 
    -- CP-element group 1202: 	1200 
    -- CP-element group 1202: 	1201 
    -- CP-element group 1202: successors 
    -- CP-element group 1202: 	696 
    -- CP-element group 1202: 	697 
    -- CP-element group 1202: 	698 
    -- CP-element group 1202: 	699 
    -- CP-element group 1202: 	700 
    -- CP-element group 1202: 	701 
    -- CP-element group 1202: 	702 
    -- CP-element group 1202: 	703 
    -- CP-element group 1202: 	704 
    -- CP-element group 1202: 	705 
    -- CP-element group 1202: 	706 
    -- CP-element group 1202: 	707 
    -- CP-element group 1202: 	709 
    -- CP-element group 1202: 	711 
    -- CP-element group 1202: 	713 
    -- CP-element group 1202: 	715 
    -- CP-element group 1202: 	717 
    -- CP-element group 1202:  members (79) 
      -- CP-element group 1202: 	 branch_block_stmt_655/merge_stmt_4343__exit__
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460__entry__
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_sample_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_Sample/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_Sample/rr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4359_Update/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_sample_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_Sample/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_Sample/rr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4369_Update/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_sample_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_word_address_calculated
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_root_address_calculated
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Sample/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Sample/word_access_start/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Sample/word_access_start/word_0/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Sample/word_access_start/word_0/rr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/word_access_complete/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/word_access_complete/word_0/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_pad_4384_Update/word_access_complete/word_0/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_sample_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_word_address_calculated
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_root_address_calculated
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Sample/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Sample/word_access_start/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Sample/word_access_start/word_0/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Sample/word_access_start/word_0/rr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/word_access_complete/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/word_access_complete/word_0/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_depth_high_4387_Update/word_access_complete/word_0/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_sample_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_word_address_calculated
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_root_address_calculated
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Sample/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Sample/word_access_start/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Sample/word_access_start/word_0/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Sample/word_access_start/word_0/rr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/word_access_complete/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/word_access_complete/word_0/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_depth_high_4390_Update/word_access_complete/word_0/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_sample_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_word_address_calculated
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_root_address_calculated
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Sample/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Sample/word_access_start/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Sample/word_access_start/word_0/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Sample/word_access_start/word_0/rr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/word_access_complete/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/word_access_complete/word_0/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/LOAD_out_col_high_4393_Update/word_access_complete/word_0/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4397_Update/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4401_Update/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4405_Update/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4414_Update/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_update_start_
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_Update/$entry
      -- CP-element group 1202: 	 branch_block_stmt_655/assign_stmt_4360_to_assign_stmt_4460/type_cast_4418_Update/cr
      -- CP-element group 1202: 	 branch_block_stmt_655/merge_stmt_4343_PhiAck/$exit
      -- 
    rr_9629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4359_inst_req_0); -- 
    cr_9634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4359_inst_req_1); -- 
    rr_9643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4369_inst_req_0); -- 
    cr_9648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4369_inst_req_1); -- 
    rr_9665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => LOAD_pad_4384_load_0_req_0); -- 
    cr_9676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => LOAD_pad_4384_load_0_req_1); -- 
    rr_9698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => LOAD_depth_high_4387_load_0_req_0); -- 
    cr_9709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => LOAD_depth_high_4387_load_0_req_1); -- 
    rr_9731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => LOAD_out_depth_high_4390_load_0_req_0); -- 
    cr_9742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => LOAD_out_depth_high_4390_load_0_req_1); -- 
    rr_9764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => LOAD_out_col_high_4393_load_0_req_0); -- 
    cr_9775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => LOAD_out_col_high_4393_load_0_req_1); -- 
    cr_9794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4397_inst_req_1); -- 
    cr_9808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4401_inst_req_1); -- 
    cr_9822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4405_inst_req_1); -- 
    cr_9836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4414_inst_req_1); -- 
    cr_9850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1202), ack => type_cast_4418_inst_req_1); -- 
    zeropad3D_cp_element_group_1202: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1202"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1199) & zeropad3D_CP_2067_elements(1200) & zeropad3D_CP_2067_elements(1201);
      gj_zeropad3D_cp_element_group_1202 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1203:  transition  input  bypass 
    -- CP-element group 1203: predecessors 
    -- CP-element group 1203: 	8 
    -- CP-element group 1203: successors 
    -- CP-element group 1203: 	1205 
    -- CP-element group 1203:  members (2) 
      -- CP-element group 1203: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/Sample/$exit
      -- CP-element group 1203: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/Sample/ra
      -- 
    ra_13644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4469_inst_ack_0, ack => zeropad3D_CP_2067_elements(1203)); -- 
    -- CP-element group 1204:  transition  input  bypass 
    -- CP-element group 1204: predecessors 
    -- CP-element group 1204: 	8 
    -- CP-element group 1204: successors 
    -- CP-element group 1204: 	1205 
    -- CP-element group 1204:  members (2) 
      -- CP-element group 1204: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/Update/$exit
      -- CP-element group 1204: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/Update/ca
      -- 
    ca_13649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4469_inst_ack_1, ack => zeropad3D_CP_2067_elements(1204)); -- 
    -- CP-element group 1205:  join  transition  output  bypass 
    -- CP-element group 1205: predecessors 
    -- CP-element group 1205: 	1203 
    -- CP-element group 1205: 	1204 
    -- CP-element group 1205: successors 
    -- CP-element group 1205: 	1212 
    -- CP-element group 1205:  members (5) 
      -- CP-element group 1205: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/$exit
      -- CP-element group 1205: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/$exit
      -- CP-element group 1205: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/$exit
      -- CP-element group 1205: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4469/SplitProtocol/$exit
      -- CP-element group 1205: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_req
      -- 
    phi_stmt_4463_req_13650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4463_req_13650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1205), ack => phi_stmt_4463_req_1); -- 
    zeropad3D_cp_element_group_1205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1203) & zeropad3D_CP_2067_elements(1204);
      gj_zeropad3D_cp_element_group_1205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1206:  transition  input  bypass 
    -- CP-element group 1206: predecessors 
    -- CP-element group 1206: 	8 
    -- CP-element group 1206: successors 
    -- CP-element group 1206: 	1208 
    -- CP-element group 1206:  members (2) 
      -- CP-element group 1206: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/Sample/$exit
      -- CP-element group 1206: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/Sample/ra
      -- 
    ra_13667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4475_inst_ack_0, ack => zeropad3D_CP_2067_elements(1206)); -- 
    -- CP-element group 1207:  transition  input  bypass 
    -- CP-element group 1207: predecessors 
    -- CP-element group 1207: 	8 
    -- CP-element group 1207: successors 
    -- CP-element group 1207: 	1208 
    -- CP-element group 1207:  members (2) 
      -- CP-element group 1207: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/Update/$exit
      -- CP-element group 1207: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/Update/ca
      -- 
    ca_13672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4475_inst_ack_1, ack => zeropad3D_CP_2067_elements(1207)); -- 
    -- CP-element group 1208:  join  transition  output  bypass 
    -- CP-element group 1208: predecessors 
    -- CP-element group 1208: 	1206 
    -- CP-element group 1208: 	1207 
    -- CP-element group 1208: successors 
    -- CP-element group 1208: 	1212 
    -- CP-element group 1208:  members (5) 
      -- CP-element group 1208: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/$exit
      -- CP-element group 1208: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/$exit
      -- CP-element group 1208: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/$exit
      -- CP-element group 1208: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4475/SplitProtocol/$exit
      -- CP-element group 1208: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_req
      -- 
    phi_stmt_4470_req_13673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4470_req_13673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1208), ack => phi_stmt_4470_req_1); -- 
    zeropad3D_cp_element_group_1208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1206) & zeropad3D_CP_2067_elements(1207);
      gj_zeropad3D_cp_element_group_1208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1209:  transition  input  bypass 
    -- CP-element group 1209: predecessors 
    -- CP-element group 1209: 	8 
    -- CP-element group 1209: successors 
    -- CP-element group 1209: 	1211 
    -- CP-element group 1209:  members (2) 
      -- CP-element group 1209: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/Sample/$exit
      -- CP-element group 1209: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/Sample/ra
      -- 
    ra_13690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4481_inst_ack_0, ack => zeropad3D_CP_2067_elements(1209)); -- 
    -- CP-element group 1210:  transition  input  bypass 
    -- CP-element group 1210: predecessors 
    -- CP-element group 1210: 	8 
    -- CP-element group 1210: successors 
    -- CP-element group 1210: 	1211 
    -- CP-element group 1210:  members (2) 
      -- CP-element group 1210: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/Update/$exit
      -- CP-element group 1210: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/Update/ca
      -- 
    ca_13695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4481_inst_ack_1, ack => zeropad3D_CP_2067_elements(1210)); -- 
    -- CP-element group 1211:  join  transition  output  bypass 
    -- CP-element group 1211: predecessors 
    -- CP-element group 1211: 	1209 
    -- CP-element group 1211: 	1210 
    -- CP-element group 1211: successors 
    -- CP-element group 1211: 	1212 
    -- CP-element group 1211:  members (5) 
      -- CP-element group 1211: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/$exit
      -- CP-element group 1211: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/$exit
      -- CP-element group 1211: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/$exit
      -- CP-element group 1211: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4481/SplitProtocol/$exit
      -- CP-element group 1211: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_req
      -- 
    phi_stmt_4476_req_13696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4476_req_13696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1211), ack => phi_stmt_4476_req_1); -- 
    zeropad3D_cp_element_group_1211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1209) & zeropad3D_CP_2067_elements(1210);
      gj_zeropad3D_cp_element_group_1211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1212:  join  transition  bypass 
    -- CP-element group 1212: predecessors 
    -- CP-element group 1212: 	1205 
    -- CP-element group 1212: 	1208 
    -- CP-element group 1212: 	1211 
    -- CP-element group 1212: successors 
    -- CP-element group 1212: 	1221 
    -- CP-element group 1212:  members (1) 
      -- CP-element group 1212: 	 branch_block_stmt_655/ifx_xend1705_whilex_xbody1552_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1212: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1212"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1205) & zeropad3D_CP_2067_elements(1208) & zeropad3D_CP_2067_elements(1211);
      gj_zeropad3D_cp_element_group_1212 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1213:  transition  output  delay-element  bypass 
    -- CP-element group 1213: predecessors 
    -- CP-element group 1213: 	718 
    -- CP-element group 1213: successors 
    -- CP-element group 1213: 	1220 
    -- CP-element group 1213:  members (4) 
      -- CP-element group 1213: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4463/$exit
      -- CP-element group 1213: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/$exit
      -- CP-element group 1213: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_sources/type_cast_4467_konst_delay_trans
      -- CP-element group 1213: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4463/phi_stmt_4463_req
      -- 
    phi_stmt_4463_req_13707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4463_req_13707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1213), ack => phi_stmt_4463_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(1213) is a control-delay.
    cp_element_1213_delay: control_delay_element  generic map(name => " 1213_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(718), ack => zeropad3D_CP_2067_elements(1213), clk => clk, reset =>reset);
    -- CP-element group 1214:  transition  input  bypass 
    -- CP-element group 1214: predecessors 
    -- CP-element group 1214: 	718 
    -- CP-element group 1214: successors 
    -- CP-element group 1214: 	1216 
    -- CP-element group 1214:  members (2) 
      -- CP-element group 1214: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/Sample/$exit
      -- CP-element group 1214: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/Sample/ra
      -- 
    ra_13724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4473_inst_ack_0, ack => zeropad3D_CP_2067_elements(1214)); -- 
    -- CP-element group 1215:  transition  input  bypass 
    -- CP-element group 1215: predecessors 
    -- CP-element group 1215: 	718 
    -- CP-element group 1215: successors 
    -- CP-element group 1215: 	1216 
    -- CP-element group 1215:  members (2) 
      -- CP-element group 1215: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/Update/$exit
      -- CP-element group 1215: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/Update/ca
      -- 
    ca_13729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4473_inst_ack_1, ack => zeropad3D_CP_2067_elements(1215)); -- 
    -- CP-element group 1216:  join  transition  output  bypass 
    -- CP-element group 1216: predecessors 
    -- CP-element group 1216: 	1214 
    -- CP-element group 1216: 	1215 
    -- CP-element group 1216: successors 
    -- CP-element group 1216: 	1220 
    -- CP-element group 1216:  members (5) 
      -- CP-element group 1216: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/$exit
      -- CP-element group 1216: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/$exit
      -- CP-element group 1216: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/$exit
      -- CP-element group 1216: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_sources/type_cast_4473/SplitProtocol/$exit
      -- CP-element group 1216: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4470/phi_stmt_4470_req
      -- 
    phi_stmt_4470_req_13730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4470_req_13730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1216), ack => phi_stmt_4470_req_0); -- 
    zeropad3D_cp_element_group_1216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1214) & zeropad3D_CP_2067_elements(1215);
      gj_zeropad3D_cp_element_group_1216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1217:  transition  input  bypass 
    -- CP-element group 1217: predecessors 
    -- CP-element group 1217: 	718 
    -- CP-element group 1217: successors 
    -- CP-element group 1217: 	1219 
    -- CP-element group 1217:  members (2) 
      -- CP-element group 1217: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/Sample/$exit
      -- CP-element group 1217: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/Sample/ra
      -- 
    ra_13747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4479_inst_ack_0, ack => zeropad3D_CP_2067_elements(1217)); -- 
    -- CP-element group 1218:  transition  input  bypass 
    -- CP-element group 1218: predecessors 
    -- CP-element group 1218: 	718 
    -- CP-element group 1218: successors 
    -- CP-element group 1218: 	1219 
    -- CP-element group 1218:  members (2) 
      -- CP-element group 1218: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/Update/$exit
      -- CP-element group 1218: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/Update/ca
      -- 
    ca_13752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4479_inst_ack_1, ack => zeropad3D_CP_2067_elements(1218)); -- 
    -- CP-element group 1219:  join  transition  output  bypass 
    -- CP-element group 1219: predecessors 
    -- CP-element group 1219: 	1217 
    -- CP-element group 1219: 	1218 
    -- CP-element group 1219: successors 
    -- CP-element group 1219: 	1220 
    -- CP-element group 1219:  members (5) 
      -- CP-element group 1219: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/$exit
      -- CP-element group 1219: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/$exit
      -- CP-element group 1219: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/$exit
      -- CP-element group 1219: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_sources/type_cast_4479/SplitProtocol/$exit
      -- CP-element group 1219: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/phi_stmt_4476/phi_stmt_4476_req
      -- 
    phi_stmt_4476_req_13753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4476_req_13753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1219), ack => phi_stmt_4476_req_0); -- 
    zeropad3D_cp_element_group_1219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1217) & zeropad3D_CP_2067_elements(1218);
      gj_zeropad3D_cp_element_group_1219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1220:  join  transition  bypass 
    -- CP-element group 1220: predecessors 
    -- CP-element group 1220: 	1213 
    -- CP-element group 1220: 	1216 
    -- CP-element group 1220: 	1219 
    -- CP-element group 1220: successors 
    -- CP-element group 1220: 	1221 
    -- CP-element group 1220:  members (1) 
      -- CP-element group 1220: 	 branch_block_stmt_655/whilex_xend1487_whilex_xbody1552_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1220: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1220"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1213) & zeropad3D_CP_2067_elements(1216) & zeropad3D_CP_2067_elements(1219);
      gj_zeropad3D_cp_element_group_1220 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1221:  merge  fork  transition  place  bypass 
    -- CP-element group 1221: predecessors 
    -- CP-element group 1221: 	1212 
    -- CP-element group 1221: 	1220 
    -- CP-element group 1221: successors 
    -- CP-element group 1221: 	1222 
    -- CP-element group 1221: 	1223 
    -- CP-element group 1221: 	1224 
    -- CP-element group 1221:  members (2) 
      -- CP-element group 1221: 	 branch_block_stmt_655/merge_stmt_4462_PhiReqMerge
      -- CP-element group 1221: 	 branch_block_stmt_655/merge_stmt_4462_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1221) <= OrReduce(zeropad3D_CP_2067_elements(1212) & zeropad3D_CP_2067_elements(1220));
    -- CP-element group 1222:  transition  input  bypass 
    -- CP-element group 1222: predecessors 
    -- CP-element group 1222: 	1221 
    -- CP-element group 1222: successors 
    -- CP-element group 1222: 	1225 
    -- CP-element group 1222:  members (1) 
      -- CP-element group 1222: 	 branch_block_stmt_655/merge_stmt_4462_PhiAck/phi_stmt_4463_ack
      -- 
    phi_stmt_4463_ack_13758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4463_ack_0, ack => zeropad3D_CP_2067_elements(1222)); -- 
    -- CP-element group 1223:  transition  input  bypass 
    -- CP-element group 1223: predecessors 
    -- CP-element group 1223: 	1221 
    -- CP-element group 1223: successors 
    -- CP-element group 1223: 	1225 
    -- CP-element group 1223:  members (1) 
      -- CP-element group 1223: 	 branch_block_stmt_655/merge_stmt_4462_PhiAck/phi_stmt_4470_ack
      -- 
    phi_stmt_4470_ack_13759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4470_ack_0, ack => zeropad3D_CP_2067_elements(1223)); -- 
    -- CP-element group 1224:  transition  input  bypass 
    -- CP-element group 1224: predecessors 
    -- CP-element group 1224: 	1221 
    -- CP-element group 1224: successors 
    -- CP-element group 1224: 	1225 
    -- CP-element group 1224:  members (1) 
      -- CP-element group 1224: 	 branch_block_stmt_655/merge_stmt_4462_PhiAck/phi_stmt_4476_ack
      -- 
    phi_stmt_4476_ack_13760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4476_ack_0, ack => zeropad3D_CP_2067_elements(1224)); -- 
    -- CP-element group 1225:  join  fork  transition  place  output  bypass 
    -- CP-element group 1225: predecessors 
    -- CP-element group 1225: 	1222 
    -- CP-element group 1225: 	1223 
    -- CP-element group 1225: 	1224 
    -- CP-element group 1225: successors 
    -- CP-element group 1225: 	719 
    -- CP-element group 1225: 	720 
    -- CP-element group 1225:  members (10) 
      -- CP-element group 1225: 	 branch_block_stmt_655/merge_stmt_4462__exit__
      -- CP-element group 1225: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494__entry__
      -- CP-element group 1225: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/$entry
      -- CP-element group 1225: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_sample_start_
      -- CP-element group 1225: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_update_start_
      -- CP-element group 1225: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_Sample/$entry
      -- CP-element group 1225: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_Sample/rr
      -- CP-element group 1225: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_Update/$entry
      -- CP-element group 1225: 	 branch_block_stmt_655/assign_stmt_4487_to_assign_stmt_4494/type_cast_4486_Update/cr
      -- CP-element group 1225: 	 branch_block_stmt_655/merge_stmt_4462_PhiAck/$exit
      -- 
    rr_9862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1225), ack => type_cast_4486_inst_req_0); -- 
    cr_9867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1225), ack => type_cast_4486_inst_req_1); -- 
    zeropad3D_cp_element_group_1225: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1225"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1222) & zeropad3D_CP_2067_elements(1223) & zeropad3D_CP_2067_elements(1224);
      gj_zeropad3D_cp_element_group_1225 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1226:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1226: predecessors 
    -- CP-element group 1226: 	721 
    -- CP-element group 1226: 	728 
    -- CP-element group 1226: 	731 
    -- CP-element group 1226: 	738 
    -- CP-element group 1226: successors 
    -- CP-element group 1226: 	739 
    -- CP-element group 1226: 	740 
    -- CP-element group 1226: 	741 
    -- CP-element group 1226: 	742 
    -- CP-element group 1226: 	745 
    -- CP-element group 1226: 	747 
    -- CP-element group 1226: 	749 
    -- CP-element group 1226: 	751 
    -- CP-element group 1226:  members (33) 
      -- CP-element group 1226: 	 branch_block_stmt_655/merge_stmt_4572__exit__
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628__entry__
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_sample_start_
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_update_start_
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Update/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_Update/cr
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_Update/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_Sample/rr
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_Sample/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_update_start_
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4581_sample_start_
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_Update/cr
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_Update/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_Sample/rr
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Update/word_access_complete/word_0/cr
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_Sample/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4576_update_start_
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_update_start_
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_update_start_
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_complete/req
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_Update/cr
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/addr_of_4622_complete/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_Update/req
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/type_cast_4615_Update/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_Update/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Update/word_access_complete/word_0/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/ptr_deref_4625_Update/word_access_complete/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/assign_stmt_4577_to_assign_stmt_4628/array_obj_ref_4621_final_index_sum_regn_update_start
      -- CP-element group 1226: 	 branch_block_stmt_655/merge_stmt_4572_PhiReqMerge
      -- CP-element group 1226: 	 branch_block_stmt_655/merge_stmt_4572_PhiAck/$entry
      -- CP-element group 1226: 	 branch_block_stmt_655/merge_stmt_4572_PhiAck/$exit
      -- CP-element group 1226: 	 branch_block_stmt_655/merge_stmt_4572_PhiAck/dummy
      -- 
    cr_10091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1226), ack => type_cast_4581_inst_req_1); -- 
    rr_10086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1226), ack => type_cast_4581_inst_req_0); -- 
    cr_10077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1226), ack => type_cast_4576_inst_req_1); -- 
    rr_10072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1226), ack => type_cast_4576_inst_req_0); -- 
    cr_10201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1226), ack => ptr_deref_4625_store_0_req_1); -- 
    req_10151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1226), ack => addr_of_4622_final_reg_req_1); -- 
    cr_10105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1226), ack => type_cast_4615_inst_req_1); -- 
    req_10136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1226), ack => array_obj_ref_4621_index_offset_req_1); -- 
    zeropad3D_CP_2067_elements(1226) <= OrReduce(zeropad3D_CP_2067_elements(721) & zeropad3D_CP_2067_elements(728) & zeropad3D_CP_2067_elements(731) & zeropad3D_CP_2067_elements(738));
    -- CP-element group 1227:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1227: predecessors 
    -- CP-element group 1227: 	752 
    -- CP-element group 1227: 	772 
    -- CP-element group 1227: successors 
    -- CP-element group 1227: 	773 
    -- CP-element group 1227: 	774 
    -- CP-element group 1227:  members (13) 
      -- CP-element group 1227: 	 branch_block_stmt_655/merge_stmt_4737__exit__
      -- CP-element group 1227: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755__entry__
      -- CP-element group 1227: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/$entry
      -- CP-element group 1227: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_sample_start_
      -- CP-element group 1227: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_update_start_
      -- CP-element group 1227: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_Sample/$entry
      -- CP-element group 1227: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_Sample/rr
      -- CP-element group 1227: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_Update/$entry
      -- CP-element group 1227: 	 branch_block_stmt_655/assign_stmt_4742_to_assign_stmt_4755/type_cast_4741_Update/cr
      -- CP-element group 1227: 	 branch_block_stmt_655/merge_stmt_4737_PhiReqMerge
      -- CP-element group 1227: 	 branch_block_stmt_655/merge_stmt_4737_PhiAck/$entry
      -- CP-element group 1227: 	 branch_block_stmt_655/merge_stmt_4737_PhiAck/$exit
      -- CP-element group 1227: 	 branch_block_stmt_655/merge_stmt_4737_PhiAck/dummy
      -- 
    rr_10450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1227), ack => type_cast_4741_inst_req_0); -- 
    cr_10455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1227), ack => type_cast_4741_inst_req_1); -- 
    zeropad3D_CP_2067_elements(1227) <= OrReduce(zeropad3D_CP_2067_elements(752) & zeropad3D_CP_2067_elements(772));
    -- CP-element group 1228:  transition  input  bypass 
    -- CP-element group 1228: predecessors 
    -- CP-element group 1228: 	794 
    -- CP-element group 1228: successors 
    -- CP-element group 1228: 	1230 
    -- CP-element group 1228:  members (2) 
      -- CP-element group 1228: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/Sample/$exit
      -- CP-element group 1228: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/Sample/ra
      -- 
    ra_13880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4861_inst_ack_0, ack => zeropad3D_CP_2067_elements(1228)); -- 
    -- CP-element group 1229:  transition  input  bypass 
    -- CP-element group 1229: predecessors 
    -- CP-element group 1229: 	794 
    -- CP-element group 1229: successors 
    -- CP-element group 1229: 	1230 
    -- CP-element group 1229:  members (2) 
      -- CP-element group 1229: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/Update/$exit
      -- CP-element group 1229: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/Update/ca
      -- 
    ca_13885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4861_inst_ack_1, ack => zeropad3D_CP_2067_elements(1229)); -- 
    -- CP-element group 1230:  join  transition  output  bypass 
    -- CP-element group 1230: predecessors 
    -- CP-element group 1230: 	1228 
    -- CP-element group 1230: 	1229 
    -- CP-element group 1230: successors 
    -- CP-element group 1230: 	1235 
    -- CP-element group 1230:  members (5) 
      -- CP-element group 1230: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/$exit
      -- CP-element group 1230: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/$exit
      -- CP-element group 1230: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/$exit
      -- CP-element group 1230: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4861/SplitProtocol/$exit
      -- CP-element group 1230: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_req
      -- 
    phi_stmt_4856_req_13886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4856_req_13886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1230), ack => phi_stmt_4856_req_1); -- 
    zeropad3D_cp_element_group_1230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1228) & zeropad3D_CP_2067_elements(1229);
      gj_zeropad3D_cp_element_group_1230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1231:  transition  output  delay-element  bypass 
    -- CP-element group 1231: predecessors 
    -- CP-element group 1231: 	794 
    -- CP-element group 1231: successors 
    -- CP-element group 1231: 	1235 
    -- CP-element group 1231:  members (4) 
      -- CP-element group 1231: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4843/$exit
      -- CP-element group 1231: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/$exit
      -- CP-element group 1231: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4847_konst_delay_trans
      -- CP-element group 1231: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_req
      -- 
    phi_stmt_4843_req_13894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4843_req_13894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1231), ack => phi_stmt_4843_req_0); -- 
    -- Element group zeropad3D_CP_2067_elements(1231) is a control-delay.
    cp_element_1231_delay: control_delay_element  generic map(name => " 1231_delay", delay_value => 1)  port map(req => zeropad3D_CP_2067_elements(794), ack => zeropad3D_CP_2067_elements(1231), clk => clk, reset =>reset);
    -- CP-element group 1232:  transition  input  bypass 
    -- CP-element group 1232: predecessors 
    -- CP-element group 1232: 	794 
    -- CP-element group 1232: successors 
    -- CP-element group 1232: 	1234 
    -- CP-element group 1232:  members (2) 
      -- CP-element group 1232: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/Sample/$exit
      -- CP-element group 1232: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/Sample/ra
      -- 
    ra_13911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4855_inst_ack_0, ack => zeropad3D_CP_2067_elements(1232)); -- 
    -- CP-element group 1233:  transition  input  bypass 
    -- CP-element group 1233: predecessors 
    -- CP-element group 1233: 	794 
    -- CP-element group 1233: successors 
    -- CP-element group 1233: 	1234 
    -- CP-element group 1233:  members (2) 
      -- CP-element group 1233: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/Update/$exit
      -- CP-element group 1233: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/Update/ca
      -- 
    ca_13916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4855_inst_ack_1, ack => zeropad3D_CP_2067_elements(1233)); -- 
    -- CP-element group 1234:  join  transition  output  bypass 
    -- CP-element group 1234: predecessors 
    -- CP-element group 1234: 	1232 
    -- CP-element group 1234: 	1233 
    -- CP-element group 1234: successors 
    -- CP-element group 1234: 	1235 
    -- CP-element group 1234:  members (5) 
      -- CP-element group 1234: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/$exit
      -- CP-element group 1234: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/$exit
      -- CP-element group 1234: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/$exit
      -- CP-element group 1234: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4855/SplitProtocol/$exit
      -- CP-element group 1234: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_req
      -- 
    phi_stmt_4850_req_13917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4850_req_13917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1234), ack => phi_stmt_4850_req_1); -- 
    zeropad3D_cp_element_group_1234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1232) & zeropad3D_CP_2067_elements(1233);
      gj_zeropad3D_cp_element_group_1234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1235:  join  transition  bypass 
    -- CP-element group 1235: predecessors 
    -- CP-element group 1235: 	1230 
    -- CP-element group 1235: 	1231 
    -- CP-element group 1235: 	1234 
    -- CP-element group 1235: successors 
    -- CP-element group 1235: 	1246 
    -- CP-element group 1235:  members (1) 
      -- CP-element group 1235: 	 branch_block_stmt_655/ifx_xelse1670_ifx_xend1705_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1235: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1235"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1230) & zeropad3D_CP_2067_elements(1231) & zeropad3D_CP_2067_elements(1234);
      gj_zeropad3D_cp_element_group_1235 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1236:  transition  input  bypass 
    -- CP-element group 1236: predecessors 
    -- CP-element group 1236: 	775 
    -- CP-element group 1236: successors 
    -- CP-element group 1236: 	1238 
    -- CP-element group 1236:  members (2) 
      -- CP-element group 1236: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/Sample/$exit
      -- CP-element group 1236: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/Sample/ra
      -- 
    ra_13937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4859_inst_ack_0, ack => zeropad3D_CP_2067_elements(1236)); -- 
    -- CP-element group 1237:  transition  input  bypass 
    -- CP-element group 1237: predecessors 
    -- CP-element group 1237: 	775 
    -- CP-element group 1237: successors 
    -- CP-element group 1237: 	1238 
    -- CP-element group 1237:  members (2) 
      -- CP-element group 1237: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/Update/$exit
      -- CP-element group 1237: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/Update/ca
      -- 
    ca_13942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4859_inst_ack_1, ack => zeropad3D_CP_2067_elements(1237)); -- 
    -- CP-element group 1238:  join  transition  output  bypass 
    -- CP-element group 1238: predecessors 
    -- CP-element group 1238: 	1236 
    -- CP-element group 1238: 	1237 
    -- CP-element group 1238: successors 
    -- CP-element group 1238: 	1245 
    -- CP-element group 1238:  members (5) 
      -- CP-element group 1238: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/$exit
      -- CP-element group 1238: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/$exit
      -- CP-element group 1238: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/$exit
      -- CP-element group 1238: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_sources/type_cast_4859/SplitProtocol/$exit
      -- CP-element group 1238: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4856/phi_stmt_4856_req
      -- 
    phi_stmt_4856_req_13943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4856_req_13943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1238), ack => phi_stmt_4856_req_0); -- 
    zeropad3D_cp_element_group_1238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1236) & zeropad3D_CP_2067_elements(1237);
      gj_zeropad3D_cp_element_group_1238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1239:  transition  input  bypass 
    -- CP-element group 1239: predecessors 
    -- CP-element group 1239: 	775 
    -- CP-element group 1239: successors 
    -- CP-element group 1239: 	1241 
    -- CP-element group 1239:  members (2) 
      -- CP-element group 1239: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/Sample/$exit
      -- CP-element group 1239: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/Sample/ra
      -- 
    ra_13960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4849_inst_ack_0, ack => zeropad3D_CP_2067_elements(1239)); -- 
    -- CP-element group 1240:  transition  input  bypass 
    -- CP-element group 1240: predecessors 
    -- CP-element group 1240: 	775 
    -- CP-element group 1240: successors 
    -- CP-element group 1240: 	1241 
    -- CP-element group 1240:  members (2) 
      -- CP-element group 1240: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/Update/$exit
      -- CP-element group 1240: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/Update/ca
      -- 
    ca_13965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4849_inst_ack_1, ack => zeropad3D_CP_2067_elements(1240)); -- 
    -- CP-element group 1241:  join  transition  output  bypass 
    -- CP-element group 1241: predecessors 
    -- CP-element group 1241: 	1239 
    -- CP-element group 1241: 	1240 
    -- CP-element group 1241: successors 
    -- CP-element group 1241: 	1245 
    -- CP-element group 1241:  members (5) 
      -- CP-element group 1241: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/$exit
      -- CP-element group 1241: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/$exit
      -- CP-element group 1241: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/$exit
      -- CP-element group 1241: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_sources/type_cast_4849/SplitProtocol/$exit
      -- CP-element group 1241: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4843/phi_stmt_4843_req
      -- 
    phi_stmt_4843_req_13966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4843_req_13966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1241), ack => phi_stmt_4843_req_1); -- 
    zeropad3D_cp_element_group_1241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1239) & zeropad3D_CP_2067_elements(1240);
      gj_zeropad3D_cp_element_group_1241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1242:  transition  input  bypass 
    -- CP-element group 1242: predecessors 
    -- CP-element group 1242: 	775 
    -- CP-element group 1242: successors 
    -- CP-element group 1242: 	1244 
    -- CP-element group 1242:  members (2) 
      -- CP-element group 1242: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/Sample/$exit
      -- CP-element group 1242: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/Sample/ra
      -- 
    ra_13983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4853_inst_ack_0, ack => zeropad3D_CP_2067_elements(1242)); -- 
    -- CP-element group 1243:  transition  input  bypass 
    -- CP-element group 1243: predecessors 
    -- CP-element group 1243: 	775 
    -- CP-element group 1243: successors 
    -- CP-element group 1243: 	1244 
    -- CP-element group 1243:  members (2) 
      -- CP-element group 1243: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/Update/$exit
      -- CP-element group 1243: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/Update/ca
      -- 
    ca_13988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4853_inst_ack_1, ack => zeropad3D_CP_2067_elements(1243)); -- 
    -- CP-element group 1244:  join  transition  output  bypass 
    -- CP-element group 1244: predecessors 
    -- CP-element group 1244: 	1242 
    -- CP-element group 1244: 	1243 
    -- CP-element group 1244: successors 
    -- CP-element group 1244: 	1245 
    -- CP-element group 1244:  members (5) 
      -- CP-element group 1244: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/$exit
      -- CP-element group 1244: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/$exit
      -- CP-element group 1244: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/$exit
      -- CP-element group 1244: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_sources/type_cast_4853/SplitProtocol/$exit
      -- CP-element group 1244: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/phi_stmt_4850/phi_stmt_4850_req
      -- 
    phi_stmt_4850_req_13989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4850_req_13989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2067_elements(1244), ack => phi_stmt_4850_req_0); -- 
    zeropad3D_cp_element_group_1244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1242) & zeropad3D_CP_2067_elements(1243);
      gj_zeropad3D_cp_element_group_1244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1245:  join  transition  bypass 
    -- CP-element group 1245: predecessors 
    -- CP-element group 1245: 	1238 
    -- CP-element group 1245: 	1241 
    -- CP-element group 1245: 	1244 
    -- CP-element group 1245: successors 
    -- CP-element group 1245: 	1246 
    -- CP-element group 1245:  members (1) 
      -- CP-element group 1245: 	 branch_block_stmt_655/ifx_xthen1665_ifx_xend1705_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1238) & zeropad3D_CP_2067_elements(1241) & zeropad3D_CP_2067_elements(1244);
      gj_zeropad3D_cp_element_group_1245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1246:  merge  fork  transition  place  bypass 
    -- CP-element group 1246: predecessors 
    -- CP-element group 1246: 	1235 
    -- CP-element group 1246: 	1245 
    -- CP-element group 1246: successors 
    -- CP-element group 1246: 	1247 
    -- CP-element group 1246: 	1248 
    -- CP-element group 1246: 	1249 
    -- CP-element group 1246:  members (2) 
      -- CP-element group 1246: 	 branch_block_stmt_655/merge_stmt_4842_PhiReqMerge
      -- CP-element group 1246: 	 branch_block_stmt_655/merge_stmt_4842_PhiAck/$entry
      -- 
    zeropad3D_CP_2067_elements(1246) <= OrReduce(zeropad3D_CP_2067_elements(1235) & zeropad3D_CP_2067_elements(1245));
    -- CP-element group 1247:  transition  input  bypass 
    -- CP-element group 1247: predecessors 
    -- CP-element group 1247: 	1246 
    -- CP-element group 1247: successors 
    -- CP-element group 1247: 	1250 
    -- CP-element group 1247:  members (1) 
      -- CP-element group 1247: 	 branch_block_stmt_655/merge_stmt_4842_PhiAck/phi_stmt_4843_ack
      -- 
    phi_stmt_4843_ack_13994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4843_ack_0, ack => zeropad3D_CP_2067_elements(1247)); -- 
    -- CP-element group 1248:  transition  input  bypass 
    -- CP-element group 1248: predecessors 
    -- CP-element group 1248: 	1246 
    -- CP-element group 1248: successors 
    -- CP-element group 1248: 	1250 
    -- CP-element group 1248:  members (1) 
      -- CP-element group 1248: 	 branch_block_stmt_655/merge_stmt_4842_PhiAck/phi_stmt_4850_ack
      -- 
    phi_stmt_4850_ack_13995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4850_ack_0, ack => zeropad3D_CP_2067_elements(1248)); -- 
    -- CP-element group 1249:  transition  input  bypass 
    -- CP-element group 1249: predecessors 
    -- CP-element group 1249: 	1246 
    -- CP-element group 1249: successors 
    -- CP-element group 1249: 	1250 
    -- CP-element group 1249:  members (1) 
      -- CP-element group 1249: 	 branch_block_stmt_655/merge_stmt_4842_PhiAck/phi_stmt_4856_ack
      -- 
    phi_stmt_4856_ack_13996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4856_ack_0, ack => zeropad3D_CP_2067_elements(1249)); -- 
    -- CP-element group 1250:  join  transition  bypass 
    -- CP-element group 1250: predecessors 
    -- CP-element group 1250: 	1247 
    -- CP-element group 1250: 	1248 
    -- CP-element group 1250: 	1249 
    -- CP-element group 1250: successors 
    -- CP-element group 1250: 	8 
    -- CP-element group 1250:  members (1) 
      -- CP-element group 1250: 	 branch_block_stmt_655/merge_stmt_4842_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1250: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1250"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2067_elements(1247) & zeropad3D_CP_2067_elements(1248) & zeropad3D_CP_2067_elements(1249);
      gj_zeropad3D_cp_element_group_1250 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2067_elements(1250), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1016_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1245_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1271_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1429_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1512_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1537_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1759_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1785_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1949_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2032_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2057_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2300_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2326_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2483_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2566_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2591_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2813_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2839_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3009_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3092_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3117_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3366_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3392_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3555_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3638_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3663_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3897_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3923_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4081_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4164_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4189_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4432_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4458_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4609_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4692_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4717_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_716_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_742_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_907_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_991_wire : std_logic_vector(31 downto 0);
    signal LOAD_col_high_1082_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1082_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1368_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1368_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1603_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1603_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1882_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1882_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2123_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2123_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2422_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2422_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2657_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2657_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2942_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2942_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3183_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3183_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3494_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3494_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3729_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3729_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4014_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4014_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4255_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4255_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4548_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4548_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4783_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4783_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_666_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_666_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_840_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_840_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_1200_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_1200_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_1714_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_1714_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_2255_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_2255_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_2768_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_2768_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_3321_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_3321_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_3852_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_3852_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_4387_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_4387_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_663_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_663_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_col_high_1206_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_1206_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_col_high_1720_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_1720_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_col_high_2261_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_2261_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_col_high_2774_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_2774_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_col_high_3327_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_3327_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_col_high_3858_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_3858_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_col_high_4393_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_4393_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_col_high_672_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_col_high_672_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_1203_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_1203_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_1717_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_1717_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_2258_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_2258_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_2771_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_2771_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_3324_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_3324_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_3855_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_3855_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_4390_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_4390_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_out_depth_high_669_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_out_depth_high_669_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_1197_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1197_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_1711_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1711_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_2252_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_2252_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_2765_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_2765_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_3318_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_3318_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_3849_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_3849_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_4384_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_4384_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_660_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_660_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1126_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1126_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1317_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1317_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1640_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1640_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1831_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1831_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2167_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2167_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2371_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2371_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2694_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2694_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2885_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2885_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3227_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3227_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3437_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3437_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3766_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3766_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3969_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3969_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4299_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4299_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4503_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4503_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4820_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4820_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_789_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_789_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom1167_3566_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1167_3566_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom120_1002_resized : std_logic_vector(13 downto 0);
    signal R_idxprom120_1002_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1210_3649_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1210_3649_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1215_3674_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1215_3674_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom125_1027_resized : std_logic_vector(13 downto 0);
    signal R_idxprom125_1027_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1385_4092_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1385_4092_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1428_4175_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1428_4175_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1433_4200_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1433_4200_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1605_4620_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1605_4620_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1648_4703_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1648_4703_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1653_4728_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1653_4728_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom288_1440_resized : std_logic_vector(13 downto 0);
    signal R_idxprom288_1440_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom331_1523_resized : std_logic_vector(13 downto 0);
    signal R_idxprom331_1523_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom336_1548_resized : std_logic_vector(13 downto 0);
    signal R_idxprom336_1548_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom505_1960_resized : std_logic_vector(13 downto 0);
    signal R_idxprom505_1960_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom548_2043_resized : std_logic_vector(13 downto 0);
    signal R_idxprom548_2043_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom553_2068_resized : std_logic_vector(13 downto 0);
    signal R_idxprom553_2068_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom726_2494_resized : std_logic_vector(13 downto 0);
    signal R_idxprom726_2494_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom769_2577_resized : std_logic_vector(13 downto 0);
    signal R_idxprom769_2577_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom774_2602_resized : std_logic_vector(13 downto 0);
    signal R_idxprom774_2602_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom944_3020_resized : std_logic_vector(13 downto 0);
    signal R_idxprom944_3020_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom987_3103_resized : std_logic_vector(13 downto 0);
    signal R_idxprom987_3103_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom992_3128_resized : std_logic_vector(13 downto 0);
    signal R_idxprom992_3128_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_919_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_919_scaled : std_logic_vector(13 downto 0);
    signal add1007_3168 : std_logic_vector(15 downto 0);
    signal add101_964 : std_logic_vector(31 downto 0);
    signal add1020_3199 : std_logic_vector(31 downto 0);
    signal add1037_3249 : std_logic_vector(31 downto 0);
    signal add111_979 : std_logic_vector(31 downto 0);
    signal add1128_3459 : std_logic_vector(31 downto 0);
    signal add1145_3504 : std_logic_vector(31 downto 0);
    signal add1158_3543 : std_logic_vector(31 downto 0);
    signal add1164_3548 : std_logic_vector(31 downto 0);
    signal add117_984 : std_logic_vector(31 downto 0);
    signal add1182_3606 : std_logic_vector(31 downto 0);
    signal add1191_3611 : std_logic_vector(31 downto 0);
    signal add1201_3626 : std_logic_vector(31 downto 0);
    signal add1207_3631 : std_logic_vector(31 downto 0);
    signal add1222_3694 : std_logic_vector(31 downto 0);
    signal add1230_3714 : std_logic_vector(15 downto 0);
    signal add1242_3739 : std_logic_vector(31 downto 0);
    signal add1259_3788 : std_logic_vector(31 downto 0);
    signal add130_1047 : std_logic_vector(31 downto 0);
    signal add1345_3979 : std_logic_vector(31 downto 0);
    signal add1363_4030 : std_logic_vector(31 downto 0);
    signal add1376_4069 : std_logic_vector(31 downto 0);
    signal add1382_4074 : std_logic_vector(31 downto 0);
    signal add138_1067 : std_logic_vector(15 downto 0);
    signal add1400_4132 : std_logic_vector(31 downto 0);
    signal add1409_4137 : std_logic_vector(31 downto 0);
    signal add1419_4152 : std_logic_vector(31 downto 0);
    signal add1425_4157 : std_logic_vector(31 downto 0);
    signal add1440_4220 : std_logic_vector(31 downto 0);
    signal add1448_4240 : std_logic_vector(15 downto 0);
    signal add1461_4271 : std_logic_vector(31 downto 0);
    signal add1476_4309 : std_logic_vector(31 downto 0);
    signal add149_1098 : std_logic_vector(31 downto 0);
    signal add1566_4513 : std_logic_vector(31 downto 0);
    signal add1583_4558 : std_logic_vector(31 downto 0);
    signal add1596_4597 : std_logic_vector(31 downto 0);
    signal add1602_4602 : std_logic_vector(31 downto 0);
    signal add1620_4660 : std_logic_vector(31 downto 0);
    signal add1629_4665 : std_logic_vector(31 downto 0);
    signal add1639_4680 : std_logic_vector(31 downto 0);
    signal add1645_4685 : std_logic_vector(31 downto 0);
    signal add165_1142 : std_logic_vector(31 downto 0);
    signal add1660_4748 : std_logic_vector(31 downto 0);
    signal add1668_4768 : std_logic_vector(15 downto 0);
    signal add1680_4793 : std_logic_vector(31 downto 0);
    signal add1695_4830 : std_logic_vector(31 downto 0);
    signal add249_1333 : std_logic_vector(31 downto 0);
    signal add266_1378 : std_logic_vector(31 downto 0);
    signal add279_1417 : std_logic_vector(31 downto 0);
    signal add285_1422 : std_logic_vector(31 downto 0);
    signal add303_1480 : std_logic_vector(31 downto 0);
    signal add312_1485 : std_logic_vector(31 downto 0);
    signal add322_1500 : std_logic_vector(31 downto 0);
    signal add328_1505 : std_logic_vector(31 downto 0);
    signal add343_1568 : std_logic_vector(31 downto 0);
    signal add351_1588 : std_logic_vector(15 downto 0);
    signal add363_1613 : std_logic_vector(31 downto 0);
    signal add379_1656 : std_logic_vector(31 downto 0);
    signal add465_1847 : std_logic_vector(31 downto 0);
    signal add483_1898 : std_logic_vector(31 downto 0);
    signal add496_1937 : std_logic_vector(31 downto 0);
    signal add502_1942 : std_logic_vector(31 downto 0);
    signal add520_2000 : std_logic_vector(31 downto 0);
    signal add529_2005 : std_logic_vector(31 downto 0);
    signal add539_2020 : std_logic_vector(31 downto 0);
    signal add545_2025 : std_logic_vector(31 downto 0);
    signal add560_2088 : std_logic_vector(31 downto 0);
    signal add568_2108 : std_logic_vector(15 downto 0);
    signal add581_2139 : std_logic_vector(31 downto 0);
    signal add597_2183 : std_logic_vector(31 downto 0);
    signal add63_856 : std_logic_vector(31 downto 0);
    signal add687_2387 : std_logic_vector(31 downto 0);
    signal add704_2432 : std_logic_vector(31 downto 0);
    signal add717_2471 : std_logic_vector(31 downto 0);
    signal add723_2476 : std_logic_vector(31 downto 0);
    signal add741_2534 : std_logic_vector(31 downto 0);
    signal add74_895 : std_logic_vector(31 downto 0);
    signal add750_2539 : std_logic_vector(31 downto 0);
    signal add760_2554 : std_logic_vector(31 downto 0);
    signal add766_2559 : std_logic_vector(31 downto 0);
    signal add781_2622 : std_logic_vector(31 downto 0);
    signal add789_2642 : std_logic_vector(15 downto 0);
    signal add801_2667 : std_logic_vector(31 downto 0);
    signal add80_900 : std_logic_vector(31 downto 0);
    signal add817_2710 : std_logic_vector(31 downto 0);
    signal add904_2907 : std_logic_vector(31 downto 0);
    signal add922_2958 : std_logic_vector(31 downto 0);
    signal add92_959 : std_logic_vector(31 downto 0);
    signal add935_2997 : std_logic_vector(31 downto 0);
    signal add941_3002 : std_logic_vector(31 downto 0);
    signal add959_3060 : std_logic_vector(31 downto 0);
    signal add968_3065 : std_logic_vector(31 downto 0);
    signal add978_3080 : std_logic_vector(31 downto 0);
    signal add984_3085 : std_logic_vector(31 downto 0);
    signal add999_3148 : std_logic_vector(31 downto 0);
    signal add_805 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1003_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1003_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1003_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1003_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1003_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1003_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1028_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1028_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1028_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1028_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1028_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1028_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1441_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1441_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1441_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1441_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1441_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1441_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2044_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2044_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2044_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2044_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2044_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2044_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2069_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2069_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2069_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2069_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2069_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2069_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2495_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2578_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2578_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2578_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2578_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2578_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2578_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2603_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2603_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2603_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2603_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2603_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2603_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3021_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3021_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3021_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3021_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3021_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3021_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3104_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3104_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3104_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3104_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3104_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3104_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3129_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3129_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3129_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3129_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3129_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3129_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3567_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3567_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3567_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3567_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3567_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3567_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3650_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3650_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3650_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3650_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3650_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3650_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3675_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3675_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3675_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3675_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3675_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3675_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4093_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4093_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4093_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4093_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4093_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4093_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4176_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4176_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4176_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4176_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4176_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4176_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4201_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4201_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4201_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4201_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4201_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4201_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4621_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4621_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4621_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4621_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4621_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4621_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4704_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4704_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4704_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4704_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4704_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4704_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4729_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4729_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4729_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4729_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4729_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4729_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_920_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_920_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_920_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_920_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_920_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_920_root_address : std_logic_vector(13 downto 0);
    signal arrayidx1168_3569 : std_logic_vector(31 downto 0);
    signal arrayidx1211_3652 : std_logic_vector(31 downto 0);
    signal arrayidx1216_3677 : std_logic_vector(31 downto 0);
    signal arrayidx121_1005 : std_logic_vector(31 downto 0);
    signal arrayidx126_1030 : std_logic_vector(31 downto 0);
    signal arrayidx1386_4095 : std_logic_vector(31 downto 0);
    signal arrayidx1429_4178 : std_logic_vector(31 downto 0);
    signal arrayidx1434_4203 : std_logic_vector(31 downto 0);
    signal arrayidx1606_4623 : std_logic_vector(31 downto 0);
    signal arrayidx1649_4706 : std_logic_vector(31 downto 0);
    signal arrayidx1654_4731 : std_logic_vector(31 downto 0);
    signal arrayidx289_1443 : std_logic_vector(31 downto 0);
    signal arrayidx332_1526 : std_logic_vector(31 downto 0);
    signal arrayidx337_1551 : std_logic_vector(31 downto 0);
    signal arrayidx506_1963 : std_logic_vector(31 downto 0);
    signal arrayidx549_2046 : std_logic_vector(31 downto 0);
    signal arrayidx554_2071 : std_logic_vector(31 downto 0);
    signal arrayidx727_2497 : std_logic_vector(31 downto 0);
    signal arrayidx770_2580 : std_logic_vector(31 downto 0);
    signal arrayidx775_2605 : std_logic_vector(31 downto 0);
    signal arrayidx945_3023 : std_logic_vector(31 downto 0);
    signal arrayidx988_3106 : std_logic_vector(31 downto 0);
    signal arrayidx993_3131 : std_logic_vector(31 downto 0);
    signal arrayidx_922 : std_logic_vector(31 downto 0);
    signal call_657 : std_logic_vector(15 downto 0);
    signal cmp1002_3155 : std_logic_vector(0 downto 0);
    signal cmp1021_3204 : std_logic_vector(0 downto 0);
    signal cmp1038_3254 : std_logic_vector(0 downto 0);
    signal cmp1117_3428 : std_logic_vector(0 downto 0);
    signal cmp1129_3466 : std_logic_vector(0 downto 0);
    signal cmp1136_3485 : std_logic_vector(0 downto 0);
    signal cmp1146_3511 : std_logic_vector(0 downto 0);
    signal cmp1225_3701 : std_logic_vector(0 downto 0);
    signal cmp1243_3744 : std_logic_vector(0 downto 0);
    signal cmp1260_3793 : std_logic_vector(0 downto 0);
    signal cmp1336_3960 : std_logic_vector(0 downto 0);
    signal cmp133_1054 : std_logic_vector(0 downto 0);
    signal cmp1346_3986 : std_logic_vector(0 downto 0);
    signal cmp1353_4005 : std_logic_vector(0 downto 0);
    signal cmp1364_4037 : std_logic_vector(0 downto 0);
    signal cmp1443_4227 : std_logic_vector(0 downto 0);
    signal cmp1462_4276 : std_logic_vector(0 downto 0);
    signal cmp1477_4314 : std_logic_vector(0 downto 0);
    signal cmp150_1103 : std_logic_vector(0 downto 0);
    signal cmp1557_4494 : std_logic_vector(0 downto 0);
    signal cmp1567_4520 : std_logic_vector(0 downto 0);
    signal cmp1574_4539 : std_logic_vector(0 downto 0);
    signal cmp1584_4565 : std_logic_vector(0 downto 0);
    signal cmp1663_4755 : std_logic_vector(0 downto 0);
    signal cmp166_1147 : std_logic_vector(0 downto 0);
    signal cmp1681_4798 : std_logic_vector(0 downto 0);
    signal cmp1696_4835 : std_logic_vector(0 downto 0);
    signal cmp239_1308 : std_logic_vector(0 downto 0);
    signal cmp250_1340 : std_logic_vector(0 downto 0);
    signal cmp257_1359 : std_logic_vector(0 downto 0);
    signal cmp267_1385 : std_logic_vector(0 downto 0);
    signal cmp346_1575 : std_logic_vector(0 downto 0);
    signal cmp364_1618 : std_logic_vector(0 downto 0);
    signal cmp380_1661 : std_logic_vector(0 downto 0);
    signal cmp455_1822 : std_logic_vector(0 downto 0);
    signal cmp466_1854 : std_logic_vector(0 downto 0);
    signal cmp46_812 : std_logic_vector(0 downto 0);
    signal cmp473_1873 : std_logic_vector(0 downto 0);
    signal cmp484_1905 : std_logic_vector(0 downto 0);
    signal cmp53_831 : std_logic_vector(0 downto 0);
    signal cmp563_2095 : std_logic_vector(0 downto 0);
    signal cmp582_2144 : std_logic_vector(0 downto 0);
    signal cmp598_2188 : std_logic_vector(0 downto 0);
    signal cmp64_863 : std_logic_vector(0 downto 0);
    signal cmp677_2362 : std_logic_vector(0 downto 0);
    signal cmp688_2394 : std_logic_vector(0 downto 0);
    signal cmp695_2413 : std_logic_vector(0 downto 0);
    signal cmp705_2439 : std_logic_vector(0 downto 0);
    signal cmp784_2629 : std_logic_vector(0 downto 0);
    signal cmp802_2672 : std_logic_vector(0 downto 0);
    signal cmp818_2715 : std_logic_vector(0 downto 0);
    signal cmp893_2876 : std_logic_vector(0 downto 0);
    signal cmp905_2914 : std_logic_vector(0 downto 0);
    signal cmp912_2933 : std_logic_vector(0 downto 0);
    signal cmp923_2965 : std_logic_vector(0 downto 0);
    signal cmp_780 : std_logic_vector(0 downto 0);
    signal conv1013_3181 : std_logic_vector(31 downto 0);
    signal conv1015_3188 : std_logic_vector(31 downto 0);
    signal conv1015x_xlcssa_3288 : std_logic_vector(31 downto 0);
    signal conv1029_3225 : std_logic_vector(31 downto 0);
    signal conv1031_3232 : std_logic_vector(31 downto 0);
    signal conv1054_3300 : std_logic_vector(15 downto 0);
    signal conv1060_3310 : std_logic_vector(15 downto 0);
    signal conv1094_3332 : std_logic_vector(31 downto 0);
    signal conv1102_3336 : std_logic_vector(31 downto 0);
    signal conv1104_3340 : std_logic_vector(31 downto 0);
    signal conv1114_3421 : std_logic_vector(31 downto 0);
    signal conv1116_3349 : std_logic_vector(31 downto 0);
    signal conv1123_3442 : std_logic_vector(31 downto 0);
    signal conv1133_3478 : std_logic_vector(31 downto 0);
    signal conv1142_3499 : std_logic_vector(31 downto 0);
    signal conv1152_3523 : std_logic_vector(31 downto 0);
    signal conv1154_3353 : std_logic_vector(31 downto 0);
    signal conv1156_3528 : std_logic_vector(31 downto 0);
    signal conv1160_3368 : std_logic_vector(31 downto 0);
    signal conv1173_3581 : std_logic_vector(31 downto 0);
    signal conv1184_3394 : std_logic_vector(31 downto 0);
    signal conv1221_3688 : std_logic_vector(31 downto 0);
    signal conv1236_3727 : std_logic_vector(31 downto 0);
    signal conv1238_3734 : std_logic_vector(31 downto 0);
    signal conv1238x_xlcssa_3827 : std_logic_vector(31 downto 0);
    signal conv1251_3764 : std_logic_vector(31 downto 0);
    signal conv1253_3771 : std_logic_vector(31 downto 0);
    signal conv1278_3835 : std_logic_vector(15 downto 0);
    signal conv129_1041 : std_logic_vector(31 downto 0);
    signal conv1313_3863 : std_logic_vector(31 downto 0);
    signal conv1321_3867 : std_logic_vector(31 downto 0);
    signal conv1323_3871 : std_logic_vector(31 downto 0);
    signal conv1333_3953 : std_logic_vector(31 downto 0);
    signal conv1335_3880 : std_logic_vector(31 downto 0);
    signal conv1342_3974 : std_logic_vector(31 downto 0);
    signal conv1350_3998 : std_logic_vector(31 downto 0);
    signal conv1359_4019 : std_logic_vector(31 downto 0);
    signal conv1370_4049 : std_logic_vector(31 downto 0);
    signal conv1372_3884 : std_logic_vector(31 downto 0);
    signal conv1374_4054 : std_logic_vector(31 downto 0);
    signal conv1378_3899 : std_logic_vector(31 downto 0);
    signal conv1391_4107 : std_logic_vector(31 downto 0);
    signal conv1402_3925 : std_logic_vector(31 downto 0);
    signal conv1439_4214 : std_logic_vector(31 downto 0);
    signal conv143_1080 : std_logic_vector(31 downto 0);
    signal conv1454_4253 : std_logic_vector(31 downto 0);
    signal conv1456_4260 : std_logic_vector(31 downto 0);
    signal conv1456x_xlcssa_4348 : std_logic_vector(31 downto 0);
    signal conv145_1087 : std_logic_vector(31 downto 0);
    signal conv145x_xlcssa_1177 : std_logic_vector(31 downto 0);
    signal conv1470_4297 : std_logic_vector(31 downto 0);
    signal conv1472_4304 : std_logic_vector(31 downto 0);
    signal conv1493_4360 : std_logic_vector(15 downto 0);
    signal conv1499_4370 : std_logic_vector(15 downto 0);
    signal conv1534_4398 : std_logic_vector(31 downto 0);
    signal conv1542_4402 : std_logic_vector(31 downto 0);
    signal conv1544_4406 : std_logic_vector(31 downto 0);
    signal conv1554_4487 : std_logic_vector(31 downto 0);
    signal conv1556_4415 : std_logic_vector(31 downto 0);
    signal conv1563_4508 : std_logic_vector(31 downto 0);
    signal conv1571_4532 : std_logic_vector(31 downto 0);
    signal conv1580_4553 : std_logic_vector(31 downto 0);
    signal conv158_1124 : std_logic_vector(31 downto 0);
    signal conv1590_4577 : std_logic_vector(31 downto 0);
    signal conv1592_4419 : std_logic_vector(31 downto 0);
    signal conv1594_4582 : std_logic_vector(31 downto 0);
    signal conv1598_4434 : std_logic_vector(31 downto 0);
    signal conv160_1131 : std_logic_vector(31 downto 0);
    signal conv1611_4635 : std_logic_vector(31 downto 0);
    signal conv1622_4460 : std_logic_vector(31 downto 0);
    signal conv1659_4742 : std_logic_vector(31 downto 0);
    signal conv1674_4781 : std_logic_vector(31 downto 0);
    signal conv1676_4788 : std_logic_vector(31 downto 0);
    signal conv1689_4818 : std_logic_vector(31 downto 0);
    signal conv1691_4825 : std_logic_vector(31 downto 0);
    signal conv180_1189 : std_logic_vector(15 downto 0);
    signal conv216_1211 : std_logic_vector(31 downto 0);
    signal conv21_677 : std_logic_vector(31 downto 0);
    signal conv224_1215 : std_logic_vector(31 downto 0);
    signal conv226_1219 : std_logic_vector(31 downto 0);
    signal conv236_1301 : std_logic_vector(31 downto 0);
    signal conv238_1228 : std_logic_vector(31 downto 0);
    signal conv23_681 : std_logic_vector(31 downto 0);
    signal conv245_1322 : std_logic_vector(31 downto 0);
    signal conv254_1352 : std_logic_vector(31 downto 0);
    signal conv263_1373 : std_logic_vector(31 downto 0);
    signal conv273_1397 : std_logic_vector(31 downto 0);
    signal conv275_1232 : std_logic_vector(31 downto 0);
    signal conv277_1402 : std_logic_vector(31 downto 0);
    signal conv27_685 : std_logic_vector(31 downto 0);
    signal conv281_1247 : std_logic_vector(31 downto 0);
    signal conv294_1455 : std_logic_vector(31 downto 0);
    signal conv29_689 : std_logic_vector(31 downto 0);
    signal conv305_1273 : std_logic_vector(31 downto 0);
    signal conv342_1562 : std_logic_vector(31 downto 0);
    signal conv357_1601 : std_logic_vector(31 downto 0);
    signal conv359_1608 : std_logic_vector(31 downto 0);
    signal conv359x_xlcssa_1695 : std_logic_vector(31 downto 0);
    signal conv36_773 : std_logic_vector(31 downto 0);
    signal conv372_1638 : std_logic_vector(31 downto 0);
    signal conv374_1645 : std_logic_vector(31 downto 0);
    signal conv38_698 : std_logic_vector(31 downto 0);
    signal conv398_1703 : std_logic_vector(15 downto 0);
    signal conv432_1725 : std_logic_vector(31 downto 0);
    signal conv43_794 : std_logic_vector(31 downto 0);
    signal conv440_1729 : std_logic_vector(31 downto 0);
    signal conv442_1733 : std_logic_vector(31 downto 0);
    signal conv452_1815 : std_logic_vector(31 downto 0);
    signal conv454_1742 : std_logic_vector(31 downto 0);
    signal conv461_1836 : std_logic_vector(31 downto 0);
    signal conv470_1866 : std_logic_vector(31 downto 0);
    signal conv479_1887 : std_logic_vector(31 downto 0);
    signal conv490_1917 : std_logic_vector(31 downto 0);
    signal conv492_1746 : std_logic_vector(31 downto 0);
    signal conv494_1922 : std_logic_vector(31 downto 0);
    signal conv498_1761 : std_logic_vector(31 downto 0);
    signal conv50_824 : std_logic_vector(31 downto 0);
    signal conv511_1975 : std_logic_vector(31 downto 0);
    signal conv522_1787 : std_logic_vector(31 downto 0);
    signal conv559_2082 : std_logic_vector(31 downto 0);
    signal conv574_2121 : std_logic_vector(31 downto 0);
    signal conv576_2128 : std_logic_vector(31 downto 0);
    signal conv576x_xlcssa_2222 : std_logic_vector(31 downto 0);
    signal conv590_2165 : std_logic_vector(31 downto 0);
    signal conv592_2172 : std_logic_vector(31 downto 0);
    signal conv59_845 : std_logic_vector(31 downto 0);
    signal conv614_2234 : std_logic_vector(15 downto 0);
    signal conv620_2244 : std_logic_vector(15 downto 0);
    signal conv654_2266 : std_logic_vector(31 downto 0);
    signal conv662_2270 : std_logic_vector(31 downto 0);
    signal conv664_2274 : std_logic_vector(31 downto 0);
    signal conv674_2355 : std_logic_vector(31 downto 0);
    signal conv676_2283 : std_logic_vector(31 downto 0);
    signal conv683_2376 : std_logic_vector(31 downto 0);
    signal conv68_875 : std_logic_vector(31 downto 0);
    signal conv692_2406 : std_logic_vector(31 downto 0);
    signal conv701_2427 : std_logic_vector(31 downto 0);
    signal conv70_702 : std_logic_vector(31 downto 0);
    signal conv711_2451 : std_logic_vector(31 downto 0);
    signal conv713_2287 : std_logic_vector(31 downto 0);
    signal conv715_2456 : std_logic_vector(31 downto 0);
    signal conv719_2302 : std_logic_vector(31 downto 0);
    signal conv72_880 : std_logic_vector(31 downto 0);
    signal conv732_2509 : std_logic_vector(31 downto 0);
    signal conv743_2328 : std_logic_vector(31 downto 0);
    signal conv76_718 : std_logic_vector(31 downto 0);
    signal conv780_2616 : std_logic_vector(31 downto 0);
    signal conv795_2655 : std_logic_vector(31 downto 0);
    signal conv797_2662 : std_logic_vector(31 downto 0);
    signal conv797x_xlcssa_2749 : std_logic_vector(31 downto 0);
    signal conv810_2692 : std_logic_vector(31 downto 0);
    signal conv812_2699 : std_logic_vector(31 downto 0);
    signal conv836_2757 : std_logic_vector(15 downto 0);
    signal conv84_934 : std_logic_vector(31 downto 0);
    signal conv870_2779 : std_logic_vector(31 downto 0);
    signal conv878_2783 : std_logic_vector(31 downto 0);
    signal conv880_2787 : std_logic_vector(31 downto 0);
    signal conv890_2869 : std_logic_vector(31 downto 0);
    signal conv892_2796 : std_logic_vector(31 downto 0);
    signal conv899_2890 : std_logic_vector(31 downto 0);
    signal conv909_2926 : std_logic_vector(31 downto 0);
    signal conv918_2947 : std_logic_vector(31 downto 0);
    signal conv929_2977 : std_logic_vector(31 downto 0);
    signal conv931_2800 : std_logic_vector(31 downto 0);
    signal conv933_2982 : std_logic_vector(31 downto 0);
    signal conv937_2815 : std_logic_vector(31 downto 0);
    signal conv94_744 : std_logic_vector(31 downto 0);
    signal conv950_3035 : std_logic_vector(31 downto 0);
    signal conv961_2841 : std_logic_vector(31 downto 0);
    signal conv998_3142 : std_logic_vector(31 downto 0);
    signal div1016_3194 : std_logic_vector(31 downto 0);
    signal div1033_3244 : std_logic_vector(31 downto 0);
    signal div1055_3306 : std_logic_vector(15 downto 0);
    signal div1061_3316 : std_logic_vector(15 downto 0);
    signal div1125_3454 : std_logic_vector(31 downto 0);
    signal div1255_3783 : std_logic_vector(31 downto 0);
    signal div1279_3841 : std_logic_vector(15 downto 0);
    signal div1360_4025 : std_logic_vector(31 downto 0);
    signal div1457_4266 : std_logic_vector(31 downto 0);
    signal div146_1093 : std_logic_vector(31 downto 0);
    signal div1494_4366 : std_logic_vector(15 downto 0);
    signal div1501_4382 : std_logic_vector(15 downto 0);
    signal div161_1137 : std_logic_vector(31 downto 0);
    signal div181_1195 : std_logic_vector(15 downto 0);
    signal div246_1328 : std_logic_vector(31 downto 0);
    signal div375_1651 : std_logic_vector(31 downto 0);
    signal div399_1709 : std_logic_vector(15 downto 0);
    signal div462_1842 : std_logic_vector(31 downto 0);
    signal div480_1893 : std_logic_vector(31 downto 0);
    signal div577_2134 : std_logic_vector(31 downto 0);
    signal div593_2178 : std_logic_vector(31 downto 0);
    signal div60_851 : std_logic_vector(31 downto 0);
    signal div615_2240 : std_logic_vector(15 downto 0);
    signal div621_2250 : std_logic_vector(15 downto 0);
    signal div684_2382 : std_logic_vector(31 downto 0);
    signal div813_2705 : std_logic_vector(31 downto 0);
    signal div837_2763 : std_logic_vector(15 downto 0);
    signal div901_2902 : std_logic_vector(31 downto 0);
    signal div919_2953 : std_logic_vector(31 downto 0);
    signal div_800 : std_logic_vector(31 downto 0);
    signal i1058x_x1x_xph_3808 : std_logic_vector(15 downto 0);
    signal i1058x_x2_3404 : std_logic_vector(15 downto 0);
    signal i1276x_x1x_xph_4329 : std_logic_vector(15 downto 0);
    signal i1276x_x2_3935 : std_logic_vector(15 downto 0);
    signal i1497x_x1x_xph_4850 : std_logic_vector(15 downto 0);
    signal i1497x_x2_4470 : std_logic_vector(15 downto 0);
    signal i184x_x1x_xph_1675 : std_logic_vector(15 downto 0);
    signal i184x_x2_1282 : std_logic_vector(15 downto 0);
    signal i396x_x1x_xph_2203 : std_logic_vector(15 downto 0);
    signal i396x_x2_1797 : std_logic_vector(15 downto 0);
    signal i618x_x1x_xph_2730 : std_logic_vector(15 downto 0);
    signal i618x_x2_2338 : std_logic_vector(15 downto 0);
    signal i834x_x1x_xph_3269 : std_logic_vector(15 downto 0);
    signal i834x_x2_2851 : std_logic_vector(15 downto 0);
    signal idxprom1167_3562 : std_logic_vector(63 downto 0);
    signal idxprom120_998 : std_logic_vector(63 downto 0);
    signal idxprom1210_3645 : std_logic_vector(63 downto 0);
    signal idxprom1215_3670 : std_logic_vector(63 downto 0);
    signal idxprom125_1023 : std_logic_vector(63 downto 0);
    signal idxprom1385_4088 : std_logic_vector(63 downto 0);
    signal idxprom1428_4171 : std_logic_vector(63 downto 0);
    signal idxprom1433_4196 : std_logic_vector(63 downto 0);
    signal idxprom1605_4616 : std_logic_vector(63 downto 0);
    signal idxprom1648_4699 : std_logic_vector(63 downto 0);
    signal idxprom1653_4724 : std_logic_vector(63 downto 0);
    signal idxprom288_1436 : std_logic_vector(63 downto 0);
    signal idxprom331_1519 : std_logic_vector(63 downto 0);
    signal idxprom336_1544 : std_logic_vector(63 downto 0);
    signal idxprom505_1956 : std_logic_vector(63 downto 0);
    signal idxprom548_2039 : std_logic_vector(63 downto 0);
    signal idxprom553_2064 : std_logic_vector(63 downto 0);
    signal idxprom726_2490 : std_logic_vector(63 downto 0);
    signal idxprom769_2573 : std_logic_vector(63 downto 0);
    signal idxprom774_2598 : std_logic_vector(63 downto 0);
    signal idxprom944_3016 : std_logic_vector(63 downto 0);
    signal idxprom987_3099 : std_logic_vector(63 downto 0);
    signal idxprom992_3124 : std_logic_vector(63 downto 0);
    signal idxprom_915 : std_logic_vector(63 downto 0);
    signal inc1011_3176 : std_logic_vector(15 downto 0);
    signal inc1026_3208 : std_logic_vector(15 downto 0);
    signal inc1026x_xi834x_x2_3213 : std_logic_vector(15 downto 0);
    signal inc1234_3722 : std_logic_vector(15 downto 0);
    signal inc1248_3748 : std_logic_vector(15 downto 0);
    signal inc1248x_xi1058x_x2_3753 : std_logic_vector(15 downto 0);
    signal inc1452_4248 : std_logic_vector(15 downto 0);
    signal inc1467_4280 : std_logic_vector(15 downto 0);
    signal inc1467x_xi1276x_x2_4285 : std_logic_vector(15 downto 0);
    signal inc155_1107 : std_logic_vector(15 downto 0);
    signal inc155x_xix_x2_1112 : std_logic_vector(15 downto 0);
    signal inc1672_4776 : std_logic_vector(15 downto 0);
    signal inc1686_4802 : std_logic_vector(15 downto 0);
    signal inc1686x_xi1497x_x2_4807 : std_logic_vector(15 downto 0);
    signal inc355_1596 : std_logic_vector(15 downto 0);
    signal inc369_1622 : std_logic_vector(15 downto 0);
    signal inc369x_xi184x_x2_1627 : std_logic_vector(15 downto 0);
    signal inc572_2116 : std_logic_vector(15 downto 0);
    signal inc587_2148 : std_logic_vector(15 downto 0);
    signal inc587x_xi396x_x2_2153 : std_logic_vector(15 downto 0);
    signal inc793_2650 : std_logic_vector(15 downto 0);
    signal inc807_2676 : std_logic_vector(15 downto 0);
    signal inc807x_xi618x_x2_2681 : std_logic_vector(15 downto 0);
    signal inc_1075 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_1161 : std_logic_vector(15 downto 0);
    signal ix_x2_754 : std_logic_vector(15 downto 0);
    signal j1108x_x0x_xph_3814 : std_logic_vector(15 downto 0);
    signal j1108x_x1_3410 : std_logic_vector(15 downto 0);
    signal j1108x_x2_3759 : std_logic_vector(15 downto 0);
    signal j1327x_x0x_xph_4335 : std_logic_vector(15 downto 0);
    signal j1327x_x1_3941 : std_logic_vector(15 downto 0);
    signal j1327x_x2_4292 : std_logic_vector(15 downto 0);
    signal j1548x_x0x_xph_4856 : std_logic_vector(15 downto 0);
    signal j1548x_x1_4476 : std_logic_vector(15 downto 0);
    signal j1548x_x2_4813 : std_logic_vector(15 downto 0);
    signal j230x_x0x_xph_1669 : std_logic_vector(15 downto 0);
    signal j230x_x1_1276 : std_logic_vector(15 downto 0);
    signal j230x_x2_1633 : std_logic_vector(15 downto 0);
    signal j446x_x0x_xph_2209 : std_logic_vector(15 downto 0);
    signal j446x_x1_1803 : std_logic_vector(15 downto 0);
    signal j446x_x2_2160 : std_logic_vector(15 downto 0);
    signal j668x_x0x_xph_2736 : std_logic_vector(15 downto 0);
    signal j668x_x1_2344 : std_logic_vector(15 downto 0);
    signal j668x_x2_2687 : std_logic_vector(15 downto 0);
    signal j884x_x0x_xph_3275 : std_logic_vector(15 downto 0);
    signal j884x_x1_2857 : std_logic_vector(15 downto 0);
    signal j884x_x2_3220 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_1155 : std_logic_vector(15 downto 0);
    signal jx_x1_747 : std_logic_vector(15 downto 0);
    signal jx_x2_1119 : std_logic_vector(15 downto 0);
    signal k1050x_x0x_xph_3801 : std_logic_vector(15 downto 0);
    signal k1050x_x1_3397 : std_logic_vector(15 downto 0);
    signal k1272x_x0x_xph_4322 : std_logic_vector(15 downto 0);
    signal k1272x_x1_3928 : std_logic_vector(15 downto 0);
    signal k1489x_x0x_xph_4843 : std_logic_vector(15 downto 0);
    signal k1489x_x1_4463 : std_logic_vector(15 downto 0);
    signal k176x_x0x_xph_1681 : std_logic_vector(15 downto 0);
    signal k176x_x1_1289 : std_logic_vector(15 downto 0);
    signal k392x_x0x_xph_2196 : std_logic_vector(15 downto 0);
    signal k392x_x1_1790 : std_logic_vector(15 downto 0);
    signal k610x_x0x_xph_2723 : std_logic_vector(15 downto 0);
    signal k610x_x1_2331 : std_logic_vector(15 downto 0);
    signal k830x_x0x_xph_3262 : std_logic_vector(15 downto 0);
    signal k830x_x1_2844 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_1167 : std_logic_vector(15 downto 0);
    signal kx_x1_761 : std_logic_vector(15 downto 0);
    signal mul100_954 : std_logic_vector(31 downto 0);
    signal mul1032_3238 : std_logic_vector(31 downto 0);
    signal mul1097_3380 : std_logic_vector(31 downto 0);
    signal mul1105_3345 : std_logic_vector(31 downto 0);
    signal mul110_969 : std_logic_vector(31 downto 0);
    signal mul1124_3448 : std_logic_vector(31 downto 0);
    signal mul1157_3533 : std_logic_vector(31 downto 0);
    signal mul1163_3538 : std_logic_vector(31 downto 0);
    signal mul116_974 : std_logic_vector(31 downto 0);
    signal mul1181_3591 : std_logic_vector(31 downto 0);
    signal mul1190_3601 : std_logic_vector(31 downto 0);
    signal mul1200_3616 : std_logic_vector(31 downto 0);
    signal mul1206_3621 : std_logic_vector(31 downto 0);
    signal mul1254_3777 : std_logic_vector(31 downto 0);
    signal mul1280_3847 : std_logic_vector(15 downto 0);
    signal mul1316_3911 : std_logic_vector(31 downto 0);
    signal mul1324_3876 : std_logic_vector(31 downto 0);
    signal mul1375_4059 : std_logic_vector(31 downto 0);
    signal mul1381_4064 : std_logic_vector(31 downto 0);
    signal mul1399_4117 : std_logic_vector(31 downto 0);
    signal mul1408_4127 : std_logic_vector(31 downto 0);
    signal mul1418_4142 : std_logic_vector(31 downto 0);
    signal mul1424_4147 : std_logic_vector(31 downto 0);
    signal mul1500_4376 : std_logic_vector(15 downto 0);
    signal mul1537_4446 : std_logic_vector(31 downto 0);
    signal mul1545_4411 : std_logic_vector(31 downto 0);
    signal mul1595_4587 : std_logic_vector(31 downto 0);
    signal mul1601_4592 : std_logic_vector(31 downto 0);
    signal mul1619_4645 : std_logic_vector(31 downto 0);
    signal mul1628_4655 : std_logic_vector(31 downto 0);
    signal mul1638_4670 : std_logic_vector(31 downto 0);
    signal mul1644_4675 : std_logic_vector(31 downto 0);
    signal mul219_1259 : std_logic_vector(31 downto 0);
    signal mul227_1224 : std_logic_vector(31 downto 0);
    signal mul278_1407 : std_logic_vector(31 downto 0);
    signal mul284_1412 : std_logic_vector(31 downto 0);
    signal mul302_1465 : std_logic_vector(31 downto 0);
    signal mul30_694 : std_logic_vector(31 downto 0);
    signal mul311_1475 : std_logic_vector(31 downto 0);
    signal mul321_1490 : std_logic_vector(31 downto 0);
    signal mul327_1495 : std_logic_vector(31 downto 0);
    signal mul435_1773 : std_logic_vector(31 downto 0);
    signal mul443_1738 : std_logic_vector(31 downto 0);
    signal mul495_1927 : std_logic_vector(31 downto 0);
    signal mul501_1932 : std_logic_vector(31 downto 0);
    signal mul519_1985 : std_logic_vector(31 downto 0);
    signal mul528_1995 : std_logic_vector(31 downto 0);
    signal mul538_2010 : std_logic_vector(31 downto 0);
    signal mul544_2015 : std_logic_vector(31 downto 0);
    signal mul657_2314 : std_logic_vector(31 downto 0);
    signal mul665_2279 : std_logic_vector(31 downto 0);
    signal mul716_2461 : std_logic_vector(31 downto 0);
    signal mul722_2466 : std_logic_vector(31 downto 0);
    signal mul73_885 : std_logic_vector(31 downto 0);
    signal mul740_2519 : std_logic_vector(31 downto 0);
    signal mul749_2529 : std_logic_vector(31 downto 0);
    signal mul759_2544 : std_logic_vector(31 downto 0);
    signal mul765_2549 : std_logic_vector(31 downto 0);
    signal mul79_890 : std_logic_vector(31 downto 0);
    signal mul873_2827 : std_logic_vector(31 downto 0);
    signal mul881_2792 : std_logic_vector(31 downto 0);
    signal mul900_2896 : std_logic_vector(31 downto 0);
    signal mul91_944 : std_logic_vector(31 downto 0);
    signal mul934_2987 : std_logic_vector(31 downto 0);
    signal mul940_2992 : std_logic_vector(31 downto 0);
    signal mul958_3045 : std_logic_vector(31 downto 0);
    signal mul967_3055 : std_logic_vector(31 downto 0);
    signal mul977_3070 : std_logic_vector(31 downto 0);
    signal mul983_3075 : std_logic_vector(31 downto 0);
    signal mul_730 : std_logic_vector(31 downto 0);
    signal ptr_deref_1008_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1008_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1008_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1008_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1008_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1032_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1032_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1032_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1032_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1032_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1032_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1445_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1445_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1445_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1445_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1445_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1445_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1529_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1529_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1529_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1529_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1529_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1553_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1553_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1553_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1553_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1553_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1553_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1965_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1965_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1965_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1965_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1965_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1965_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2049_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2049_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2049_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2049_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2049_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2073_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2073_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2073_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2073_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2073_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2073_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2499_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2499_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2499_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2499_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2499_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2499_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2583_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2583_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2583_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2583_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2583_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2607_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2607_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2607_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2607_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2607_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2607_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3025_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3025_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3025_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3025_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3025_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3025_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3109_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3109_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3109_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3109_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3109_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3133_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3133_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3133_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3133_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3133_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3133_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3571_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3571_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3571_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3571_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3571_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3571_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3655_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3655_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3655_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3655_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3655_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3679_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3679_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3679_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3679_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3679_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3679_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4097_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4097_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4097_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4097_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4097_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4097_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4181_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4181_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4181_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4181_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4181_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4205_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4205_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4205_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4205_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4205_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4205_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4625_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4625_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4625_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4625_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4625_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4625_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4709_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4709_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4709_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4709_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4709_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4733_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4733_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4733_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4733_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4733_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4733_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_924_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_924_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_924_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_924_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_924_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_924_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext1707_1264 : std_logic_vector(31 downto 0);
    signal sext1708_1778 : std_logic_vector(31 downto 0);
    signal sext1709_2319 : std_logic_vector(31 downto 0);
    signal sext1710_2832 : std_logic_vector(31 downto 0);
    signal sext1711_3385 : std_logic_vector(31 downto 0);
    signal sext1712_3916 : std_logic_vector(31 downto 0);
    signal sext1713_4451 : std_logic_vector(31 downto 0);
    signal sext1746_708 : std_logic_vector(31 downto 0);
    signal sext1747_1238 : std_logic_vector(31 downto 0);
    signal sext1748_1752 : std_logic_vector(31 downto 0);
    signal sext1749_2293 : std_logic_vector(31 downto 0);
    signal sext1750_2806 : std_logic_vector(31 downto 0);
    signal sext1751_3359 : std_logic_vector(31 downto 0);
    signal sext1752_3890 : std_logic_vector(31 downto 0);
    signal sext1753_4425 : std_logic_vector(31 downto 0);
    signal sext_735 : std_logic_vector(31 downto 0);
    signal shl1019_2821 : std_logic_vector(31 downto 0);
    signal shl1241_3374 : std_logic_vector(31 downto 0);
    signal shl1460_3905 : std_logic_vector(31 downto 0);
    signal shl1679_4440 : std_logic_vector(31 downto 0);
    signal shl362_1253 : std_logic_vector(31 downto 0);
    signal shl580_1767 : std_logic_vector(31 downto 0);
    signal shl800_2308 : std_logic_vector(31 downto 0);
    signal shl_724 : std_logic_vector(31 downto 0);
    signal shr1166_3557 : std_logic_vector(31 downto 0);
    signal shr119_993 : std_logic_vector(31 downto 0);
    signal shr1209_3640 : std_logic_vector(31 downto 0);
    signal shr1214_3665 : std_logic_vector(31 downto 0);
    signal shr124_1018 : std_logic_vector(31 downto 0);
    signal shr1384_4083 : std_logic_vector(31 downto 0);
    signal shr1427_4166 : std_logic_vector(31 downto 0);
    signal shr1432_4191 : std_logic_vector(31 downto 0);
    signal shr1604_4611 : std_logic_vector(31 downto 0);
    signal shr1647_4694 : std_logic_vector(31 downto 0);
    signal shr1652_4719 : std_logic_vector(31 downto 0);
    signal shr287_1431 : std_logic_vector(31 downto 0);
    signal shr330_1514 : std_logic_vector(31 downto 0);
    signal shr335_1539 : std_logic_vector(31 downto 0);
    signal shr504_1951 : std_logic_vector(31 downto 0);
    signal shr547_2034 : std_logic_vector(31 downto 0);
    signal shr552_2059 : std_logic_vector(31 downto 0);
    signal shr725_2485 : std_logic_vector(31 downto 0);
    signal shr768_2568 : std_logic_vector(31 downto 0);
    signal shr773_2593 : std_logic_vector(31 downto 0);
    signal shr943_3011 : std_logic_vector(31 downto 0);
    signal shr986_3094 : std_logic_vector(31 downto 0);
    signal shr991_3119 : std_logic_vector(31 downto 0);
    signal shr_909 : std_logic_vector(31 downto 0);
    signal sub1180_3586 : std_logic_vector(31 downto 0);
    signal sub1189_3596 : std_logic_vector(31 downto 0);
    signal sub1398_4112 : std_logic_vector(31 downto 0);
    signal sub1407_4122 : std_logic_vector(31 downto 0);
    signal sub1618_4640 : std_logic_vector(31 downto 0);
    signal sub1627_4650 : std_logic_vector(31 downto 0);
    signal sub301_1460 : std_logic_vector(31 downto 0);
    signal sub310_1470 : std_logic_vector(31 downto 0);
    signal sub518_1980 : std_logic_vector(31 downto 0);
    signal sub527_1990 : std_logic_vector(31 downto 0);
    signal sub739_2514 : std_logic_vector(31 downto 0);
    signal sub748_2524 : std_logic_vector(31 downto 0);
    signal sub957_3040 : std_logic_vector(31 downto 0);
    signal sub966_3050 : std_logic_vector(31 downto 0);
    signal sub99_949 : std_logic_vector(31 downto 0);
    signal sub_939 : std_logic_vector(31 downto 0);
    signal tmp1014_3184 : std_logic_vector(7 downto 0);
    signal tmp1014x_xlcssa_3292 : std_logic_vector(7 downto 0);
    signal tmp1030_3228 : std_logic_vector(7 downto 0);
    signal tmp1030x_xlcssa_3284 : std_logic_vector(7 downto 0);
    signal tmp1065_3319 : std_logic_vector(7 downto 0);
    signal tmp1069_3322 : std_logic_vector(7 downto 0);
    signal tmp1081_3325 : std_logic_vector(7 downto 0);
    signal tmp1085_3328 : std_logic_vector(7 downto 0);
    signal tmp1122_3438 : std_logic_vector(7 downto 0);
    signal tmp1141_3495 : std_logic_vector(7 downto 0);
    signal tmp11_670 : std_logic_vector(7 downto 0);
    signal tmp1212_3656 : std_logic_vector(63 downto 0);
    signal tmp122_1009 : std_logic_vector(63 downto 0);
    signal tmp1237_3730 : std_logic_vector(7 downto 0);
    signal tmp1252_3767 : std_logic_vector(7 downto 0);
    signal tmp1252x_xlcssa_3823 : std_logic_vector(7 downto 0);
    signal tmp1284_3850 : std_logic_vector(7 downto 0);
    signal tmp1288_3853 : std_logic_vector(7 downto 0);
    signal tmp1300_3856 : std_logic_vector(7 downto 0);
    signal tmp1304_3859 : std_logic_vector(7 downto 0);
    signal tmp1341_3970 : std_logic_vector(7 downto 0);
    signal tmp1358_4015 : std_logic_vector(7 downto 0);
    signal tmp1430_4182 : std_logic_vector(63 downto 0);
    signal tmp144_1083 : std_logic_vector(7 downto 0);
    signal tmp144x_xlcssa_1181 : std_logic_vector(7 downto 0);
    signal tmp1455_4256 : std_logic_vector(7 downto 0);
    signal tmp1455x_xlcssa_4352 : std_logic_vector(7 downto 0);
    signal tmp1471_4300 : std_logic_vector(7 downto 0);
    signal tmp1471x_xlcssa_4344 : std_logic_vector(7 downto 0);
    signal tmp14_673 : std_logic_vector(7 downto 0);
    signal tmp1505_4385 : std_logic_vector(7 downto 0);
    signal tmp1509_4388 : std_logic_vector(7 downto 0);
    signal tmp1521_4391 : std_logic_vector(7 downto 0);
    signal tmp1525_4394 : std_logic_vector(7 downto 0);
    signal tmp1562_4504 : std_logic_vector(7 downto 0);
    signal tmp1579_4549 : std_logic_vector(7 downto 0);
    signal tmp159_1127 : std_logic_vector(7 downto 0);
    signal tmp1650_4710 : std_logic_vector(63 downto 0);
    signal tmp1675_4784 : std_logic_vector(7 downto 0);
    signal tmp1690_4821 : std_logic_vector(7 downto 0);
    signal tmp187_1198 : std_logic_vector(7 downto 0);
    signal tmp191_1201 : std_logic_vector(7 downto 0);
    signal tmp203_1204 : std_logic_vector(7 downto 0);
    signal tmp207_1207 : std_logic_vector(7 downto 0);
    signal tmp244_1318 : std_logic_vector(7 downto 0);
    signal tmp262_1369 : std_logic_vector(7 downto 0);
    signal tmp2_664 : std_logic_vector(7 downto 0);
    signal tmp333_1530 : std_logic_vector(63 downto 0);
    signal tmp358_1604 : std_logic_vector(7 downto 0);
    signal tmp373_1641 : std_logic_vector(7 downto 0);
    signal tmp373x_xlcssa_1691 : std_logic_vector(7 downto 0);
    signal tmp403_1712 : std_logic_vector(7 downto 0);
    signal tmp407_1715 : std_logic_vector(7 downto 0);
    signal tmp419_1718 : std_logic_vector(7 downto 0);
    signal tmp423_1721 : std_logic_vector(7 downto 0);
    signal tmp42_790 : std_logic_vector(7 downto 0);
    signal tmp460_1832 : std_logic_vector(7 downto 0);
    signal tmp478_1883 : std_logic_vector(7 downto 0);
    signal tmp550_2050 : std_logic_vector(63 downto 0);
    signal tmp575_2124 : std_logic_vector(7 downto 0);
    signal tmp575x_xlcssa_2226 : std_logic_vector(7 downto 0);
    signal tmp58_841 : std_logic_vector(7 downto 0);
    signal tmp591_2168 : std_logic_vector(7 downto 0);
    signal tmp591x_xlcssa_2218 : std_logic_vector(7 downto 0);
    signal tmp5_667 : std_logic_vector(7 downto 0);
    signal tmp625_2253 : std_logic_vector(7 downto 0);
    signal tmp629_2256 : std_logic_vector(7 downto 0);
    signal tmp641_2259 : std_logic_vector(7 downto 0);
    signal tmp645_2262 : std_logic_vector(7 downto 0);
    signal tmp682_2372 : std_logic_vector(7 downto 0);
    signal tmp700_2423 : std_logic_vector(7 downto 0);
    signal tmp771_2584 : std_logic_vector(63 downto 0);
    signal tmp796_2658 : std_logic_vector(7 downto 0);
    signal tmp811_2695 : std_logic_vector(7 downto 0);
    signal tmp811x_xlcssa_2745 : std_logic_vector(7 downto 0);
    signal tmp841_2766 : std_logic_vector(7 downto 0);
    signal tmp845_2769 : std_logic_vector(7 downto 0);
    signal tmp857_2772 : std_logic_vector(7 downto 0);
    signal tmp861_2775 : std_logic_vector(7 downto 0);
    signal tmp898_2886 : std_logic_vector(7 downto 0);
    signal tmp917_2943 : std_logic_vector(7 downto 0);
    signal tmp989_3110 : std_logic_vector(63 downto 0);
    signal tmp_661 : std_logic_vector(7 downto 0);
    signal type_cast_1012_wire : std_logic_vector(31 downto 0);
    signal type_cast_1015_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1021_wire : std_logic_vector(63 downto 0);
    signal type_cast_1039_wire : std_logic_vector(31 downto 0);
    signal type_cast_1045_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1050_wire : std_logic_vector(31 downto 0);
    signal type_cast_1052_wire : std_logic_vector(31 downto 0);
    signal type_cast_1065_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1073_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1078_wire : std_logic_vector(31 downto 0);
    signal type_cast_1091_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1116_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1122_wire : std_logic_vector(31 downto 0);
    signal type_cast_1135_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1158_wire : std_logic_vector(15 downto 0);
    signal type_cast_1160_wire : std_logic_vector(15 downto 0);
    signal type_cast_1164_wire : std_logic_vector(15 downto 0);
    signal type_cast_1166_wire : std_logic_vector(15 downto 0);
    signal type_cast_1170_wire : std_logic_vector(15 downto 0);
    signal type_cast_1173_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1180_wire : std_logic_vector(31 downto 0);
    signal type_cast_1184_wire : std_logic_vector(7 downto 0);
    signal type_cast_1193_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1241_wire : std_logic_vector(31 downto 0);
    signal type_cast_1244_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1251_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1257_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1267_wire : std_logic_vector(31 downto 0);
    signal type_cast_1270_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1279_wire : std_logic_vector(15 downto 0);
    signal type_cast_1281_wire : std_logic_vector(15 downto 0);
    signal type_cast_1286_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1288_wire : std_logic_vector(15 downto 0);
    signal type_cast_1293_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1295_wire : std_logic_vector(15 downto 0);
    signal type_cast_1299_wire : std_logic_vector(31 downto 0);
    signal type_cast_1304_wire : std_logic_vector(31 downto 0);
    signal type_cast_1306_wire : std_logic_vector(31 downto 0);
    signal type_cast_1326_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1336_wire : std_logic_vector(31 downto 0);
    signal type_cast_1338_wire : std_logic_vector(31 downto 0);
    signal type_cast_1350_wire : std_logic_vector(31 downto 0);
    signal type_cast_1355_wire : std_logic_vector(31 downto 0);
    signal type_cast_1357_wire : std_logic_vector(31 downto 0);
    signal type_cast_1381_wire : std_logic_vector(31 downto 0);
    signal type_cast_1383_wire : std_logic_vector(31 downto 0);
    signal type_cast_1395_wire : std_logic_vector(31 downto 0);
    signal type_cast_1400_wire : std_logic_vector(31 downto 0);
    signal type_cast_1425_wire : std_logic_vector(31 downto 0);
    signal type_cast_1428_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1434_wire : std_logic_vector(63 downto 0);
    signal type_cast_1447_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1453_wire : std_logic_vector(31 downto 0);
    signal type_cast_1508_wire : std_logic_vector(31 downto 0);
    signal type_cast_1511_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1517_wire : std_logic_vector(63 downto 0);
    signal type_cast_1533_wire : std_logic_vector(31 downto 0);
    signal type_cast_1536_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1542_wire : std_logic_vector(63 downto 0);
    signal type_cast_1560_wire : std_logic_vector(31 downto 0);
    signal type_cast_1566_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1571_wire : std_logic_vector(31 downto 0);
    signal type_cast_1573_wire : std_logic_vector(31 downto 0);
    signal type_cast_1586_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1594_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1599_wire : std_logic_vector(31 downto 0);
    signal type_cast_1636_wire : std_logic_vector(31 downto 0);
    signal type_cast_1649_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1672_wire : std_logic_vector(15 downto 0);
    signal type_cast_1674_wire : std_logic_vector(15 downto 0);
    signal type_cast_1678_wire : std_logic_vector(15 downto 0);
    signal type_cast_1680_wire : std_logic_vector(15 downto 0);
    signal type_cast_1684_wire : std_logic_vector(15 downto 0);
    signal type_cast_1687_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1694_wire : std_logic_vector(7 downto 0);
    signal type_cast_1698_wire : std_logic_vector(31 downto 0);
    signal type_cast_1707_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1750_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1755_wire : std_logic_vector(31 downto 0);
    signal type_cast_1758_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1765_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1771_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1781_wire : std_logic_vector(31 downto 0);
    signal type_cast_1784_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1793_wire : std_logic_vector(15 downto 0);
    signal type_cast_1796_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1800_wire : std_logic_vector(15 downto 0);
    signal type_cast_1802_wire : std_logic_vector(15 downto 0);
    signal type_cast_1807_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1809_wire : std_logic_vector(15 downto 0);
    signal type_cast_1813_wire : std_logic_vector(31 downto 0);
    signal type_cast_1818_wire : std_logic_vector(31 downto 0);
    signal type_cast_1820_wire : std_logic_vector(31 downto 0);
    signal type_cast_1840_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1850_wire : std_logic_vector(31 downto 0);
    signal type_cast_1852_wire : std_logic_vector(31 downto 0);
    signal type_cast_1864_wire : std_logic_vector(31 downto 0);
    signal type_cast_1869_wire : std_logic_vector(31 downto 0);
    signal type_cast_1871_wire : std_logic_vector(31 downto 0);
    signal type_cast_1891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1901_wire : std_logic_vector(31 downto 0);
    signal type_cast_1903_wire : std_logic_vector(31 downto 0);
    signal type_cast_1915_wire : std_logic_vector(31 downto 0);
    signal type_cast_1920_wire : std_logic_vector(31 downto 0);
    signal type_cast_1945_wire : std_logic_vector(31 downto 0);
    signal type_cast_1948_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1954_wire : std_logic_vector(63 downto 0);
    signal type_cast_1967_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1973_wire : std_logic_vector(31 downto 0);
    signal type_cast_2028_wire : std_logic_vector(31 downto 0);
    signal type_cast_2031_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2037_wire : std_logic_vector(63 downto 0);
    signal type_cast_2053_wire : std_logic_vector(31 downto 0);
    signal type_cast_2056_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2062_wire : std_logic_vector(63 downto 0);
    signal type_cast_2080_wire : std_logic_vector(31 downto 0);
    signal type_cast_2086_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2091_wire : std_logic_vector(31 downto 0);
    signal type_cast_2093_wire : std_logic_vector(31 downto 0);
    signal type_cast_2106_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2114_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2119_wire : std_logic_vector(31 downto 0);
    signal type_cast_2132_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2157_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2163_wire : std_logic_vector(31 downto 0);
    signal type_cast_2176_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2199_wire : std_logic_vector(15 downto 0);
    signal type_cast_2202_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2206_wire : std_logic_vector(15 downto 0);
    signal type_cast_2208_wire : std_logic_vector(15 downto 0);
    signal type_cast_2212_wire : std_logic_vector(15 downto 0);
    signal type_cast_2214_wire : std_logic_vector(15 downto 0);
    signal type_cast_2221_wire : std_logic_vector(7 downto 0);
    signal type_cast_2225_wire : std_logic_vector(31 downto 0);
    signal type_cast_2229_wire : std_logic_vector(7 downto 0);
    signal type_cast_2238_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2248_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2291_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2296_wire : std_logic_vector(31 downto 0);
    signal type_cast_2299_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2306_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2312_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2322_wire : std_logic_vector(31 downto 0);
    signal type_cast_2325_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2335_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2337_wire : std_logic_vector(15 downto 0);
    signal type_cast_2341_wire : std_logic_vector(15 downto 0);
    signal type_cast_2343_wire : std_logic_vector(15 downto 0);
    signal type_cast_2347_wire : std_logic_vector(15 downto 0);
    signal type_cast_2349_wire : std_logic_vector(15 downto 0);
    signal type_cast_2353_wire : std_logic_vector(31 downto 0);
    signal type_cast_2358_wire : std_logic_vector(31 downto 0);
    signal type_cast_2360_wire : std_logic_vector(31 downto 0);
    signal type_cast_2380_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2390_wire : std_logic_vector(31 downto 0);
    signal type_cast_2392_wire : std_logic_vector(31 downto 0);
    signal type_cast_2404_wire : std_logic_vector(31 downto 0);
    signal type_cast_2409_wire : std_logic_vector(31 downto 0);
    signal type_cast_2411_wire : std_logic_vector(31 downto 0);
    signal type_cast_2435_wire : std_logic_vector(31 downto 0);
    signal type_cast_2437_wire : std_logic_vector(31 downto 0);
    signal type_cast_2449_wire : std_logic_vector(31 downto 0);
    signal type_cast_2454_wire : std_logic_vector(31 downto 0);
    signal type_cast_2479_wire : std_logic_vector(31 downto 0);
    signal type_cast_2482_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2488_wire : std_logic_vector(63 downto 0);
    signal type_cast_2501_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2507_wire : std_logic_vector(31 downto 0);
    signal type_cast_2562_wire : std_logic_vector(31 downto 0);
    signal type_cast_2565_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2571_wire : std_logic_vector(63 downto 0);
    signal type_cast_2587_wire : std_logic_vector(31 downto 0);
    signal type_cast_2590_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2596_wire : std_logic_vector(63 downto 0);
    signal type_cast_2614_wire : std_logic_vector(31 downto 0);
    signal type_cast_2620_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2625_wire : std_logic_vector(31 downto 0);
    signal type_cast_2627_wire : std_logic_vector(31 downto 0);
    signal type_cast_2640_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2648_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2653_wire : std_logic_vector(31 downto 0);
    signal type_cast_2690_wire : std_logic_vector(31 downto 0);
    signal type_cast_2703_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2726_wire : std_logic_vector(15 downto 0);
    signal type_cast_2729_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2733_wire : std_logic_vector(15 downto 0);
    signal type_cast_2735_wire : std_logic_vector(15 downto 0);
    signal type_cast_2739_wire : std_logic_vector(15 downto 0);
    signal type_cast_2741_wire : std_logic_vector(15 downto 0);
    signal type_cast_2748_wire : std_logic_vector(7 downto 0);
    signal type_cast_2752_wire : std_logic_vector(31 downto 0);
    signal type_cast_2761_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2804_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2809_wire : std_logic_vector(31 downto 0);
    signal type_cast_2812_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2819_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2825_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2835_wire : std_logic_vector(31 downto 0);
    signal type_cast_2838_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2848_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2850_wire : std_logic_vector(15 downto 0);
    signal type_cast_2854_wire : std_logic_vector(15 downto 0);
    signal type_cast_2856_wire : std_logic_vector(15 downto 0);
    signal type_cast_2861_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2863_wire : std_logic_vector(15 downto 0);
    signal type_cast_2867_wire : std_logic_vector(31 downto 0);
    signal type_cast_2872_wire : std_logic_vector(31 downto 0);
    signal type_cast_2874_wire : std_logic_vector(31 downto 0);
    signal type_cast_2894_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2900_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2910_wire : std_logic_vector(31 downto 0);
    signal type_cast_2912_wire : std_logic_vector(31 downto 0);
    signal type_cast_2924_wire : std_logic_vector(31 downto 0);
    signal type_cast_2929_wire : std_logic_vector(31 downto 0);
    signal type_cast_2931_wire : std_logic_vector(31 downto 0);
    signal type_cast_2951_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2961_wire : std_logic_vector(31 downto 0);
    signal type_cast_2963_wire : std_logic_vector(31 downto 0);
    signal type_cast_2975_wire : std_logic_vector(31 downto 0);
    signal type_cast_2980_wire : std_logic_vector(31 downto 0);
    signal type_cast_3005_wire : std_logic_vector(31 downto 0);
    signal type_cast_3008_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3014_wire : std_logic_vector(63 downto 0);
    signal type_cast_3027_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3033_wire : std_logic_vector(31 downto 0);
    signal type_cast_3088_wire : std_logic_vector(31 downto 0);
    signal type_cast_3091_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3097_wire : std_logic_vector(63 downto 0);
    signal type_cast_3113_wire : std_logic_vector(31 downto 0);
    signal type_cast_3116_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3122_wire : std_logic_vector(63 downto 0);
    signal type_cast_3140_wire : std_logic_vector(31 downto 0);
    signal type_cast_3146_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3151_wire : std_logic_vector(31 downto 0);
    signal type_cast_3153_wire : std_logic_vector(31 downto 0);
    signal type_cast_3166_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3174_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3179_wire : std_logic_vector(31 downto 0);
    signal type_cast_3192_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3217_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3223_wire : std_logic_vector(31 downto 0);
    signal type_cast_3236_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3242_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3266_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3268_wire : std_logic_vector(15 downto 0);
    signal type_cast_3272_wire : std_logic_vector(15 downto 0);
    signal type_cast_3274_wire : std_logic_vector(15 downto 0);
    signal type_cast_3278_wire : std_logic_vector(15 downto 0);
    signal type_cast_3280_wire : std_logic_vector(15 downto 0);
    signal type_cast_3287_wire : std_logic_vector(7 downto 0);
    signal type_cast_3291_wire : std_logic_vector(31 downto 0);
    signal type_cast_3295_wire : std_logic_vector(7 downto 0);
    signal type_cast_3304_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3314_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3357_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3362_wire : std_logic_vector(31 downto 0);
    signal type_cast_3365_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3372_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3378_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3388_wire : std_logic_vector(31 downto 0);
    signal type_cast_3391_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3401_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3403_wire : std_logic_vector(15 downto 0);
    signal type_cast_3407_wire : std_logic_vector(15 downto 0);
    signal type_cast_3409_wire : std_logic_vector(15 downto 0);
    signal type_cast_3413_wire : std_logic_vector(15 downto 0);
    signal type_cast_3415_wire : std_logic_vector(15 downto 0);
    signal type_cast_3419_wire : std_logic_vector(31 downto 0);
    signal type_cast_3424_wire : std_logic_vector(31 downto 0);
    signal type_cast_3426_wire : std_logic_vector(31 downto 0);
    signal type_cast_3446_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3452_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3462_wire : std_logic_vector(31 downto 0);
    signal type_cast_3464_wire : std_logic_vector(31 downto 0);
    signal type_cast_3476_wire : std_logic_vector(31 downto 0);
    signal type_cast_3481_wire : std_logic_vector(31 downto 0);
    signal type_cast_3483_wire : std_logic_vector(31 downto 0);
    signal type_cast_3507_wire : std_logic_vector(31 downto 0);
    signal type_cast_3509_wire : std_logic_vector(31 downto 0);
    signal type_cast_3521_wire : std_logic_vector(31 downto 0);
    signal type_cast_3526_wire : std_logic_vector(31 downto 0);
    signal type_cast_3551_wire : std_logic_vector(31 downto 0);
    signal type_cast_3554_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3560_wire : std_logic_vector(63 downto 0);
    signal type_cast_3573_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3579_wire : std_logic_vector(31 downto 0);
    signal type_cast_3634_wire : std_logic_vector(31 downto 0);
    signal type_cast_3637_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3643_wire : std_logic_vector(63 downto 0);
    signal type_cast_3659_wire : std_logic_vector(31 downto 0);
    signal type_cast_3662_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3668_wire : std_logic_vector(63 downto 0);
    signal type_cast_3686_wire : std_logic_vector(31 downto 0);
    signal type_cast_3692_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3697_wire : std_logic_vector(31 downto 0);
    signal type_cast_3699_wire : std_logic_vector(31 downto 0);
    signal type_cast_3712_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3720_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3725_wire : std_logic_vector(31 downto 0);
    signal type_cast_3762_wire : std_logic_vector(31 downto 0);
    signal type_cast_3775_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3781_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3804_wire : std_logic_vector(15 downto 0);
    signal type_cast_3807_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3811_wire : std_logic_vector(15 downto 0);
    signal type_cast_3813_wire : std_logic_vector(15 downto 0);
    signal type_cast_3817_wire : std_logic_vector(15 downto 0);
    signal type_cast_3819_wire : std_logic_vector(15 downto 0);
    signal type_cast_3826_wire : std_logic_vector(7 downto 0);
    signal type_cast_3830_wire : std_logic_vector(31 downto 0);
    signal type_cast_3839_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3845_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3888_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3893_wire : std_logic_vector(31 downto 0);
    signal type_cast_3896_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3903_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3909_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3919_wire : std_logic_vector(31 downto 0);
    signal type_cast_3922_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3932_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3934_wire : std_logic_vector(15 downto 0);
    signal type_cast_3938_wire : std_logic_vector(15 downto 0);
    signal type_cast_3940_wire : std_logic_vector(15 downto 0);
    signal type_cast_3945_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3947_wire : std_logic_vector(15 downto 0);
    signal type_cast_3951_wire : std_logic_vector(31 downto 0);
    signal type_cast_3956_wire : std_logic_vector(31 downto 0);
    signal type_cast_3958_wire : std_logic_vector(31 downto 0);
    signal type_cast_3982_wire : std_logic_vector(31 downto 0);
    signal type_cast_3984_wire : std_logic_vector(31 downto 0);
    signal type_cast_3996_wire : std_logic_vector(31 downto 0);
    signal type_cast_4001_wire : std_logic_vector(31 downto 0);
    signal type_cast_4003_wire : std_logic_vector(31 downto 0);
    signal type_cast_4023_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4033_wire : std_logic_vector(31 downto 0);
    signal type_cast_4035_wire : std_logic_vector(31 downto 0);
    signal type_cast_4047_wire : std_logic_vector(31 downto 0);
    signal type_cast_4052_wire : std_logic_vector(31 downto 0);
    signal type_cast_4077_wire : std_logic_vector(31 downto 0);
    signal type_cast_4080_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4086_wire : std_logic_vector(63 downto 0);
    signal type_cast_4099_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_4105_wire : std_logic_vector(31 downto 0);
    signal type_cast_4160_wire : std_logic_vector(31 downto 0);
    signal type_cast_4163_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4169_wire : std_logic_vector(63 downto 0);
    signal type_cast_4185_wire : std_logic_vector(31 downto 0);
    signal type_cast_4188_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4194_wire : std_logic_vector(63 downto 0);
    signal type_cast_4212_wire : std_logic_vector(31 downto 0);
    signal type_cast_4218_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4223_wire : std_logic_vector(31 downto 0);
    signal type_cast_4225_wire : std_logic_vector(31 downto 0);
    signal type_cast_4238_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4246_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4251_wire : std_logic_vector(31 downto 0);
    signal type_cast_4264_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4289_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4295_wire : std_logic_vector(31 downto 0);
    signal type_cast_4325_wire : std_logic_vector(15 downto 0);
    signal type_cast_4328_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4332_wire : std_logic_vector(15 downto 0);
    signal type_cast_4334_wire : std_logic_vector(15 downto 0);
    signal type_cast_4338_wire : std_logic_vector(15 downto 0);
    signal type_cast_4340_wire : std_logic_vector(15 downto 0);
    signal type_cast_4347_wire : std_logic_vector(7 downto 0);
    signal type_cast_4351_wire : std_logic_vector(31 downto 0);
    signal type_cast_4355_wire : std_logic_vector(7 downto 0);
    signal type_cast_4364_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4374_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4380_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4423_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4428_wire : std_logic_vector(31 downto 0);
    signal type_cast_4431_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4438_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4444_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4454_wire : std_logic_vector(31 downto 0);
    signal type_cast_4457_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4467_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4469_wire : std_logic_vector(15 downto 0);
    signal type_cast_4473_wire : std_logic_vector(15 downto 0);
    signal type_cast_4475_wire : std_logic_vector(15 downto 0);
    signal type_cast_4479_wire : std_logic_vector(15 downto 0);
    signal type_cast_4481_wire : std_logic_vector(15 downto 0);
    signal type_cast_4485_wire : std_logic_vector(31 downto 0);
    signal type_cast_4490_wire : std_logic_vector(31 downto 0);
    signal type_cast_4492_wire : std_logic_vector(31 downto 0);
    signal type_cast_4516_wire : std_logic_vector(31 downto 0);
    signal type_cast_4518_wire : std_logic_vector(31 downto 0);
    signal type_cast_4530_wire : std_logic_vector(31 downto 0);
    signal type_cast_4535_wire : std_logic_vector(31 downto 0);
    signal type_cast_4537_wire : std_logic_vector(31 downto 0);
    signal type_cast_4561_wire : std_logic_vector(31 downto 0);
    signal type_cast_4563_wire : std_logic_vector(31 downto 0);
    signal type_cast_4575_wire : std_logic_vector(31 downto 0);
    signal type_cast_4580_wire : std_logic_vector(31 downto 0);
    signal type_cast_4605_wire : std_logic_vector(31 downto 0);
    signal type_cast_4608_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4614_wire : std_logic_vector(63 downto 0);
    signal type_cast_4627_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_4633_wire : std_logic_vector(31 downto 0);
    signal type_cast_4688_wire : std_logic_vector(31 downto 0);
    signal type_cast_4691_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4697_wire : std_logic_vector(63 downto 0);
    signal type_cast_4713_wire : std_logic_vector(31 downto 0);
    signal type_cast_4716_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4722_wire : std_logic_vector(63 downto 0);
    signal type_cast_4740_wire : std_logic_vector(31 downto 0);
    signal type_cast_4746_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4751_wire : std_logic_vector(31 downto 0);
    signal type_cast_4753_wire : std_logic_vector(31 downto 0);
    signal type_cast_4766_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4774_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4779_wire : std_logic_vector(31 downto 0);
    signal type_cast_4816_wire : std_logic_vector(31 downto 0);
    signal type_cast_4847_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4849_wire : std_logic_vector(15 downto 0);
    signal type_cast_4853_wire : std_logic_vector(15 downto 0);
    signal type_cast_4855_wire : std_logic_vector(15 downto 0);
    signal type_cast_4859_wire : std_logic_vector(15 downto 0);
    signal type_cast_4861_wire : std_logic_vector(15 downto 0);
    signal type_cast_706_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_712_wire : std_logic_vector(31 downto 0);
    signal type_cast_715_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_722_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_728_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_738_wire : std_logic_vector(31 downto 0);
    signal type_cast_741_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_751_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_753_wire : std_logic_vector(15 downto 0);
    signal type_cast_758_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_760_wire : std_logic_vector(15 downto 0);
    signal type_cast_765_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_767_wire : std_logic_vector(15 downto 0);
    signal type_cast_771_wire : std_logic_vector(31 downto 0);
    signal type_cast_776_wire : std_logic_vector(31 downto 0);
    signal type_cast_778_wire : std_logic_vector(31 downto 0);
    signal type_cast_798_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_808_wire : std_logic_vector(31 downto 0);
    signal type_cast_810_wire : std_logic_vector(31 downto 0);
    signal type_cast_822_wire : std_logic_vector(31 downto 0);
    signal type_cast_827_wire : std_logic_vector(31 downto 0);
    signal type_cast_829_wire : std_logic_vector(31 downto 0);
    signal type_cast_849_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_859_wire : std_logic_vector(31 downto 0);
    signal type_cast_861_wire : std_logic_vector(31 downto 0);
    signal type_cast_873_wire : std_logic_vector(31 downto 0);
    signal type_cast_878_wire : std_logic_vector(31 downto 0);
    signal type_cast_903_wire : std_logic_vector(31 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_913_wire : std_logic_vector(63 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_932_wire : std_logic_vector(31 downto 0);
    signal type_cast_987_wire : std_logic_vector(31 downto 0);
    signal type_cast_990_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_996_wire : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    LOAD_col_high_1082_word_address_0 <= "0";
    LOAD_col_high_1368_word_address_0 <= "0";
    LOAD_col_high_1603_word_address_0 <= "0";
    LOAD_col_high_1882_word_address_0 <= "0";
    LOAD_col_high_2123_word_address_0 <= "0";
    LOAD_col_high_2422_word_address_0 <= "0";
    LOAD_col_high_2657_word_address_0 <= "0";
    LOAD_col_high_2942_word_address_0 <= "0";
    LOAD_col_high_3183_word_address_0 <= "0";
    LOAD_col_high_3494_word_address_0 <= "0";
    LOAD_col_high_3729_word_address_0 <= "0";
    LOAD_col_high_4014_word_address_0 <= "0";
    LOAD_col_high_4255_word_address_0 <= "0";
    LOAD_col_high_4548_word_address_0 <= "0";
    LOAD_col_high_4783_word_address_0 <= "0";
    LOAD_col_high_666_word_address_0 <= "0";
    LOAD_col_high_840_word_address_0 <= "0";
    LOAD_depth_high_1200_word_address_0 <= "0";
    LOAD_depth_high_1714_word_address_0 <= "0";
    LOAD_depth_high_2255_word_address_0 <= "0";
    LOAD_depth_high_2768_word_address_0 <= "0";
    LOAD_depth_high_3321_word_address_0 <= "0";
    LOAD_depth_high_3852_word_address_0 <= "0";
    LOAD_depth_high_4387_word_address_0 <= "0";
    LOAD_depth_high_663_word_address_0 <= "0";
    LOAD_out_col_high_1206_word_address_0 <= "0";
    LOAD_out_col_high_1720_word_address_0 <= "0";
    LOAD_out_col_high_2261_word_address_0 <= "0";
    LOAD_out_col_high_2774_word_address_0 <= "0";
    LOAD_out_col_high_3327_word_address_0 <= "0";
    LOAD_out_col_high_3858_word_address_0 <= "0";
    LOAD_out_col_high_4393_word_address_0 <= "0";
    LOAD_out_col_high_672_word_address_0 <= "0";
    LOAD_out_depth_high_1203_word_address_0 <= "0";
    LOAD_out_depth_high_1717_word_address_0 <= "0";
    LOAD_out_depth_high_2258_word_address_0 <= "0";
    LOAD_out_depth_high_2771_word_address_0 <= "0";
    LOAD_out_depth_high_3324_word_address_0 <= "0";
    LOAD_out_depth_high_3855_word_address_0 <= "0";
    LOAD_out_depth_high_4390_word_address_0 <= "0";
    LOAD_out_depth_high_669_word_address_0 <= "0";
    LOAD_pad_1197_word_address_0 <= "0";
    LOAD_pad_1711_word_address_0 <= "0";
    LOAD_pad_2252_word_address_0 <= "0";
    LOAD_pad_2765_word_address_0 <= "0";
    LOAD_pad_3318_word_address_0 <= "0";
    LOAD_pad_3849_word_address_0 <= "0";
    LOAD_pad_4384_word_address_0 <= "0";
    LOAD_pad_660_word_address_0 <= "0";
    LOAD_row_high_1126_word_address_0 <= "0";
    LOAD_row_high_1317_word_address_0 <= "0";
    LOAD_row_high_1640_word_address_0 <= "0";
    LOAD_row_high_1831_word_address_0 <= "0";
    LOAD_row_high_2167_word_address_0 <= "0";
    LOAD_row_high_2371_word_address_0 <= "0";
    LOAD_row_high_2694_word_address_0 <= "0";
    LOAD_row_high_2885_word_address_0 <= "0";
    LOAD_row_high_3227_word_address_0 <= "0";
    LOAD_row_high_3437_word_address_0 <= "0";
    LOAD_row_high_3766_word_address_0 <= "0";
    LOAD_row_high_3969_word_address_0 <= "0";
    LOAD_row_high_4299_word_address_0 <= "0";
    LOAD_row_high_4503_word_address_0 <= "0";
    LOAD_row_high_4820_word_address_0 <= "0";
    LOAD_row_high_789_word_address_0 <= "0";
    array_obj_ref_1003_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1003_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1003_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1003_resized_base_address <= "00000000000000";
    array_obj_ref_1028_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1028_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1028_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1028_resized_base_address <= "00000000000000";
    array_obj_ref_1441_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1441_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1441_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1441_resized_base_address <= "00000000000000";
    array_obj_ref_1524_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1524_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1524_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1524_resized_base_address <= "00000000000000";
    array_obj_ref_1549_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1549_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1549_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1549_resized_base_address <= "00000000000000";
    array_obj_ref_1961_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1961_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1961_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1961_resized_base_address <= "00000000000000";
    array_obj_ref_2044_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2044_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2044_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2044_resized_base_address <= "00000000000000";
    array_obj_ref_2069_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2069_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2069_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2069_resized_base_address <= "00000000000000";
    array_obj_ref_2495_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2495_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2495_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2495_resized_base_address <= "00000000000000";
    array_obj_ref_2578_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2578_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2578_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2578_resized_base_address <= "00000000000000";
    array_obj_ref_2603_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2603_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2603_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2603_resized_base_address <= "00000000000000";
    array_obj_ref_3021_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3021_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3021_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3021_resized_base_address <= "00000000000000";
    array_obj_ref_3104_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3104_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3104_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3104_resized_base_address <= "00000000000000";
    array_obj_ref_3129_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3129_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3129_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3129_resized_base_address <= "00000000000000";
    array_obj_ref_3567_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3567_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3567_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3567_resized_base_address <= "00000000000000";
    array_obj_ref_3650_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3650_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3650_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3650_resized_base_address <= "00000000000000";
    array_obj_ref_3675_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3675_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3675_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3675_resized_base_address <= "00000000000000";
    array_obj_ref_4093_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4093_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4093_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4093_resized_base_address <= "00000000000000";
    array_obj_ref_4176_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4176_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4176_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4176_resized_base_address <= "00000000000000";
    array_obj_ref_4201_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4201_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4201_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4201_resized_base_address <= "00000000000000";
    array_obj_ref_4621_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4621_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4621_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4621_resized_base_address <= "00000000000000";
    array_obj_ref_4704_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4704_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4704_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4704_resized_base_address <= "00000000000000";
    array_obj_ref_4729_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4729_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4729_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4729_resized_base_address <= "00000000000000";
    array_obj_ref_920_constant_part_of_offset <= "00000000000000";
    array_obj_ref_920_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_920_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_920_resized_base_address <= "00000000000000";
    ptr_deref_1008_word_offset_0 <= "00000000000000";
    ptr_deref_1032_word_offset_0 <= "00000000000000";
    ptr_deref_1445_word_offset_0 <= "00000000000000";
    ptr_deref_1529_word_offset_0 <= "00000000000000";
    ptr_deref_1553_word_offset_0 <= "00000000000000";
    ptr_deref_1965_word_offset_0 <= "00000000000000";
    ptr_deref_2049_word_offset_0 <= "00000000000000";
    ptr_deref_2073_word_offset_0 <= "00000000000000";
    ptr_deref_2499_word_offset_0 <= "00000000000000";
    ptr_deref_2583_word_offset_0 <= "00000000000000";
    ptr_deref_2607_word_offset_0 <= "00000000000000";
    ptr_deref_3025_word_offset_0 <= "00000000000000";
    ptr_deref_3109_word_offset_0 <= "00000000000000";
    ptr_deref_3133_word_offset_0 <= "00000000000000";
    ptr_deref_3571_word_offset_0 <= "00000000000000";
    ptr_deref_3655_word_offset_0 <= "00000000000000";
    ptr_deref_3679_word_offset_0 <= "00000000000000";
    ptr_deref_4097_word_offset_0 <= "00000000000000";
    ptr_deref_4181_word_offset_0 <= "00000000000000";
    ptr_deref_4205_word_offset_0 <= "00000000000000";
    ptr_deref_4625_word_offset_0 <= "00000000000000";
    ptr_deref_4709_word_offset_0 <= "00000000000000";
    ptr_deref_4733_word_offset_0 <= "00000000000000";
    ptr_deref_924_word_offset_0 <= "00000000000000";
    type_cast_1015_wire_constant <= "00000000000000000000000000000010";
    type_cast_1045_wire_constant <= "00000000000000000000000000000100";
    type_cast_1065_wire_constant <= "0000000000000100";
    type_cast_1073_wire_constant <= "0000000000000001";
    type_cast_1091_wire_constant <= "00000000000000000000000000000001";
    type_cast_1116_wire_constant <= "0000000000000000";
    type_cast_1135_wire_constant <= "00000000000000000000000000000010";
    type_cast_1173_wire_constant <= "0000000000000000";
    type_cast_1193_wire_constant <= "0000000000000001";
    type_cast_1236_wire_constant <= "00000000000000000000000000010000";
    type_cast_1244_wire_constant <= "00000000000000000000000000010000";
    type_cast_1251_wire_constant <= "00000000000000000000000000000001";
    type_cast_1257_wire_constant <= "00000000000000000000000000010000";
    type_cast_1270_wire_constant <= "00000000000000000000000000010000";
    type_cast_1286_wire_constant <= "0000000000000000";
    type_cast_1293_wire_constant <= "0000000000000000";
    type_cast_1326_wire_constant <= "00000000000000000000000000000010";
    type_cast_1428_wire_constant <= "00000000000000000000000000000010";
    type_cast_1447_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1511_wire_constant <= "00000000000000000000000000000010";
    type_cast_1536_wire_constant <= "00000000000000000000000000000010";
    type_cast_1566_wire_constant <= "00000000000000000000000000000100";
    type_cast_1586_wire_constant <= "0000000000000100";
    type_cast_1594_wire_constant <= "0000000000000001";
    type_cast_1649_wire_constant <= "00000000000000000000000000000010";
    type_cast_1687_wire_constant <= "0000000000000000";
    type_cast_1707_wire_constant <= "0000000000000010";
    type_cast_1750_wire_constant <= "00000000000000000000000000010000";
    type_cast_1758_wire_constant <= "00000000000000000000000000010000";
    type_cast_1765_wire_constant <= "00000000000000000000000000000001";
    type_cast_1771_wire_constant <= "00000000000000000000000000010000";
    type_cast_1784_wire_constant <= "00000000000000000000000000010000";
    type_cast_1796_wire_constant <= "0000000000000000";
    type_cast_1807_wire_constant <= "0000000000000000";
    type_cast_1840_wire_constant <= "00000000000000000000000000000001";
    type_cast_1891_wire_constant <= "00000000000000000000000000000001";
    type_cast_1948_wire_constant <= "00000000000000000000000000000010";
    type_cast_1967_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2031_wire_constant <= "00000000000000000000000000000010";
    type_cast_2056_wire_constant <= "00000000000000000000000000000010";
    type_cast_2086_wire_constant <= "00000000000000000000000000000100";
    type_cast_2106_wire_constant <= "0000000000000100";
    type_cast_2114_wire_constant <= "0000000000000001";
    type_cast_2132_wire_constant <= "00000000000000000000000000000001";
    type_cast_2157_wire_constant <= "0000000000000000";
    type_cast_2176_wire_constant <= "00000000000000000000000000000001";
    type_cast_2202_wire_constant <= "0000000000000000";
    type_cast_2238_wire_constant <= "0000000000000001";
    type_cast_2248_wire_constant <= "0000000000000010";
    type_cast_2291_wire_constant <= "00000000000000000000000000010000";
    type_cast_2299_wire_constant <= "00000000000000000000000000010000";
    type_cast_2306_wire_constant <= "00000000000000000000000000000001";
    type_cast_2312_wire_constant <= "00000000000000000000000000010000";
    type_cast_2325_wire_constant <= "00000000000000000000000000010000";
    type_cast_2335_wire_constant <= "0000000000000000";
    type_cast_2380_wire_constant <= "00000000000000000000000000000001";
    type_cast_2482_wire_constant <= "00000000000000000000000000000010";
    type_cast_2501_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2565_wire_constant <= "00000000000000000000000000000010";
    type_cast_2590_wire_constant <= "00000000000000000000000000000010";
    type_cast_2620_wire_constant <= "00000000000000000000000000000100";
    type_cast_2640_wire_constant <= "0000000000000100";
    type_cast_2648_wire_constant <= "0000000000000001";
    type_cast_2703_wire_constant <= "00000000000000000000000000000001";
    type_cast_2729_wire_constant <= "0000000000000000";
    type_cast_2761_wire_constant <= "0000000000000001";
    type_cast_2804_wire_constant <= "00000000000000000000000000010000";
    type_cast_2812_wire_constant <= "00000000000000000000000000010000";
    type_cast_2819_wire_constant <= "00000000000000000000000000000001";
    type_cast_2825_wire_constant <= "00000000000000000000000000010000";
    type_cast_2838_wire_constant <= "00000000000000000000000000010000";
    type_cast_2848_wire_constant <= "0000000000000000";
    type_cast_2861_wire_constant <= "0000000000000000";
    type_cast_2894_wire_constant <= "00000000000000000000000000000011";
    type_cast_2900_wire_constant <= "00000000000000000000000000000010";
    type_cast_2951_wire_constant <= "00000000000000000000000000000001";
    type_cast_3008_wire_constant <= "00000000000000000000000000000010";
    type_cast_3027_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3091_wire_constant <= "00000000000000000000000000000010";
    type_cast_3116_wire_constant <= "00000000000000000000000000000010";
    type_cast_3146_wire_constant <= "00000000000000000000000000000100";
    type_cast_3166_wire_constant <= "0000000000000100";
    type_cast_3174_wire_constant <= "0000000000000001";
    type_cast_3192_wire_constant <= "00000000000000000000000000000001";
    type_cast_3217_wire_constant <= "0000000000000000";
    type_cast_3236_wire_constant <= "00000000000000000000000000000011";
    type_cast_3242_wire_constant <= "00000000000000000000000000000010";
    type_cast_3266_wire_constant <= "0000000000000000";
    type_cast_3304_wire_constant <= "0000000000000001";
    type_cast_3314_wire_constant <= "0000000000000001";
    type_cast_3357_wire_constant <= "00000000000000000000000000010000";
    type_cast_3365_wire_constant <= "00000000000000000000000000010000";
    type_cast_3372_wire_constant <= "00000000000000000000000000000001";
    type_cast_3378_wire_constant <= "00000000000000000000000000010000";
    type_cast_3391_wire_constant <= "00000000000000000000000000010000";
    type_cast_3401_wire_constant <= "0000000000000000";
    type_cast_3446_wire_constant <= "00000000000000000000000000000011";
    type_cast_3452_wire_constant <= "00000000000000000000000000000010";
    type_cast_3554_wire_constant <= "00000000000000000000000000000010";
    type_cast_3573_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3637_wire_constant <= "00000000000000000000000000000010";
    type_cast_3662_wire_constant <= "00000000000000000000000000000010";
    type_cast_3692_wire_constant <= "00000000000000000000000000000100";
    type_cast_3712_wire_constant <= "0000000000000100";
    type_cast_3720_wire_constant <= "0000000000000001";
    type_cast_3775_wire_constant <= "00000000000000000000000000000011";
    type_cast_3781_wire_constant <= "00000000000000000000000000000010";
    type_cast_3807_wire_constant <= "0000000000000000";
    type_cast_3839_wire_constant <= "0000000000000010";
    type_cast_3845_wire_constant <= "0000000000000011";
    type_cast_3888_wire_constant <= "00000000000000000000000000010000";
    type_cast_3896_wire_constant <= "00000000000000000000000000010000";
    type_cast_3903_wire_constant <= "00000000000000000000000000000001";
    type_cast_3909_wire_constant <= "00000000000000000000000000010000";
    type_cast_3922_wire_constant <= "00000000000000000000000000010000";
    type_cast_3932_wire_constant <= "0000000000000000";
    type_cast_3945_wire_constant <= "0000000000000000";
    type_cast_4023_wire_constant <= "00000000000000000000000000000001";
    type_cast_4080_wire_constant <= "00000000000000000000000000000010";
    type_cast_4099_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_4163_wire_constant <= "00000000000000000000000000000010";
    type_cast_4188_wire_constant <= "00000000000000000000000000000010";
    type_cast_4218_wire_constant <= "00000000000000000000000000000100";
    type_cast_4238_wire_constant <= "0000000000000100";
    type_cast_4246_wire_constant <= "0000000000000001";
    type_cast_4264_wire_constant <= "00000000000000000000000000000001";
    type_cast_4289_wire_constant <= "0000000000000000";
    type_cast_4328_wire_constant <= "0000000000000000";
    type_cast_4364_wire_constant <= "0000000000000001";
    type_cast_4374_wire_constant <= "0000000000000011";
    type_cast_4380_wire_constant <= "0000000000000010";
    type_cast_4423_wire_constant <= "00000000000000000000000000010000";
    type_cast_4431_wire_constant <= "00000000000000000000000000010000";
    type_cast_4438_wire_constant <= "00000000000000000000000000000001";
    type_cast_4444_wire_constant <= "00000000000000000000000000010000";
    type_cast_4457_wire_constant <= "00000000000000000000000000010000";
    type_cast_4467_wire_constant <= "0000000000000000";
    type_cast_4608_wire_constant <= "00000000000000000000000000000010";
    type_cast_4627_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_4691_wire_constant <= "00000000000000000000000000000010";
    type_cast_4716_wire_constant <= "00000000000000000000000000000010";
    type_cast_4746_wire_constant <= "00000000000000000000000000000100";
    type_cast_4766_wire_constant <= "0000000000000100";
    type_cast_4774_wire_constant <= "0000000000000001";
    type_cast_4847_wire_constant <= "0000000000000000";
    type_cast_706_wire_constant <= "00000000000000000000000000010000";
    type_cast_715_wire_constant <= "00000000000000000000000000010000";
    type_cast_722_wire_constant <= "00000000000000000000000000000001";
    type_cast_728_wire_constant <= "00000000000000000000000000010000";
    type_cast_741_wire_constant <= "00000000000000000000000000010000";
    type_cast_751_wire_constant <= "0000000000000000";
    type_cast_758_wire_constant <= "0000000000000000";
    type_cast_765_wire_constant <= "0000000000000000";
    type_cast_798_wire_constant <= "00000000000000000000000000000010";
    type_cast_849_wire_constant <= "00000000000000000000000000000001";
    type_cast_906_wire_constant <= "00000000000000000000000000000010";
    type_cast_926_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_990_wire_constant <= "00000000000000000000000000000010";
    phi_stmt_1155: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1158_wire & type_cast_1160_wire;
      req <= phi_stmt_1155_req_0 & phi_stmt_1155_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1155",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1155_ack_0,
          idata => idata,
          odata => jx_x0x_xph_1155,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1155
    phi_stmt_1161: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1164_wire & type_cast_1166_wire;
      req <= phi_stmt_1161_req_0 & phi_stmt_1161_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1161",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1161_ack_0,
          idata => idata,
          odata => ix_x1x_xph_1161,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1161
    phi_stmt_1167: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1170_wire & type_cast_1173_wire_constant;
      req <= phi_stmt_1167_req_0 & phi_stmt_1167_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1167",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1167_ack_0,
          idata => idata,
          odata => kx_x0x_xph_1167,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1167
    phi_stmt_1177: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1180_wire;
      req(0) <= phi_stmt_1177_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1177",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1177_ack_0,
          idata => idata,
          odata => conv145x_xlcssa_1177,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1177
    phi_stmt_1181: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1184_wire;
      req(0) <= phi_stmt_1181_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1181",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1181_ack_0,
          idata => idata,
          odata => tmp144x_xlcssa_1181,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1181
    phi_stmt_1276: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1279_wire & type_cast_1281_wire;
      req <= phi_stmt_1276_req_0 & phi_stmt_1276_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1276",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1276_ack_0,
          idata => idata,
          odata => j230x_x1_1276,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1276
    phi_stmt_1282: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1286_wire_constant & type_cast_1288_wire;
      req <= phi_stmt_1282_req_0 & phi_stmt_1282_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1282",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1282_ack_0,
          idata => idata,
          odata => i184x_x2_1282,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1282
    phi_stmt_1289: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1293_wire_constant & type_cast_1295_wire;
      req <= phi_stmt_1289_req_0 & phi_stmt_1289_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1289",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1289_ack_0,
          idata => idata,
          odata => k176x_x1_1289,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1289
    phi_stmt_1669: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1672_wire & type_cast_1674_wire;
      req <= phi_stmt_1669_req_0 & phi_stmt_1669_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1669",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1669_ack_0,
          idata => idata,
          odata => j230x_x0x_xph_1669,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1669
    phi_stmt_1675: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1678_wire & type_cast_1680_wire;
      req <= phi_stmt_1675_req_0 & phi_stmt_1675_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1675",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1675_ack_0,
          idata => idata,
          odata => i184x_x1x_xph_1675,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1675
    phi_stmt_1681: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1684_wire & type_cast_1687_wire_constant;
      req <= phi_stmt_1681_req_0 & phi_stmt_1681_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1681",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1681_ack_0,
          idata => idata,
          odata => k176x_x0x_xph_1681,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1681
    phi_stmt_1691: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1694_wire;
      req(0) <= phi_stmt_1691_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1691",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1691_ack_0,
          idata => idata,
          odata => tmp373x_xlcssa_1691,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1691
    phi_stmt_1695: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1698_wire;
      req(0) <= phi_stmt_1695_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1695",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1695_ack_0,
          idata => idata,
          odata => conv359x_xlcssa_1695,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1695
    phi_stmt_1790: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1793_wire & type_cast_1796_wire_constant;
      req <= phi_stmt_1790_req_0 & phi_stmt_1790_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1790",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1790_ack_0,
          idata => idata,
          odata => k392x_x1_1790,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1790
    phi_stmt_1797: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1800_wire & type_cast_1802_wire;
      req <= phi_stmt_1797_req_0 & phi_stmt_1797_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1797",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1797_ack_0,
          idata => idata,
          odata => i396x_x2_1797,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1797
    phi_stmt_1803: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1807_wire_constant & type_cast_1809_wire;
      req <= phi_stmt_1803_req_0 & phi_stmt_1803_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1803",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1803_ack_0,
          idata => idata,
          odata => j446x_x1_1803,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1803
    phi_stmt_2196: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2199_wire & type_cast_2202_wire_constant;
      req <= phi_stmt_2196_req_0 & phi_stmt_2196_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2196",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2196_ack_0,
          idata => idata,
          odata => k392x_x0x_xph_2196,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2196
    phi_stmt_2203: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2206_wire & type_cast_2208_wire;
      req <= phi_stmt_2203_req_0 & phi_stmt_2203_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2203",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2203_ack_0,
          idata => idata,
          odata => i396x_x1x_xph_2203,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2203
    phi_stmt_2209: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2212_wire & type_cast_2214_wire;
      req <= phi_stmt_2209_req_0 & phi_stmt_2209_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2209",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2209_ack_0,
          idata => idata,
          odata => j446x_x0x_xph_2209,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2209
    phi_stmt_2218: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2221_wire;
      req(0) <= phi_stmt_2218_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2218",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2218_ack_0,
          idata => idata,
          odata => tmp591x_xlcssa_2218,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2218
    phi_stmt_2222: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2225_wire;
      req(0) <= phi_stmt_2222_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2222",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2222_ack_0,
          idata => idata,
          odata => conv576x_xlcssa_2222,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2222
    phi_stmt_2226: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2229_wire;
      req(0) <= phi_stmt_2226_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2226",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2226_ack_0,
          idata => idata,
          odata => tmp575x_xlcssa_2226,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2226
    phi_stmt_2331: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2335_wire_constant & type_cast_2337_wire;
      req <= phi_stmt_2331_req_0 & phi_stmt_2331_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2331",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2331_ack_0,
          idata => idata,
          odata => k610x_x1_2331,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2331
    phi_stmt_2338: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2341_wire & type_cast_2343_wire;
      req <= phi_stmt_2338_req_0 & phi_stmt_2338_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2338",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2338_ack_0,
          idata => idata,
          odata => i618x_x2_2338,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2338
    phi_stmt_2344: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2347_wire & type_cast_2349_wire;
      req <= phi_stmt_2344_req_0 & phi_stmt_2344_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2344",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2344_ack_0,
          idata => idata,
          odata => j668x_x1_2344,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2344
    phi_stmt_2723: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2726_wire & type_cast_2729_wire_constant;
      req <= phi_stmt_2723_req_0 & phi_stmt_2723_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2723",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2723_ack_0,
          idata => idata,
          odata => k610x_x0x_xph_2723,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2723
    phi_stmt_2730: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2733_wire & type_cast_2735_wire;
      req <= phi_stmt_2730_req_0 & phi_stmt_2730_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2730",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2730_ack_0,
          idata => idata,
          odata => i618x_x1x_xph_2730,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2730
    phi_stmt_2736: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2739_wire & type_cast_2741_wire;
      req <= phi_stmt_2736_req_0 & phi_stmt_2736_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2736",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2736_ack_0,
          idata => idata,
          odata => j668x_x0x_xph_2736,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2736
    phi_stmt_2745: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2748_wire;
      req(0) <= phi_stmt_2745_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2745",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2745_ack_0,
          idata => idata,
          odata => tmp811x_xlcssa_2745,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2745
    phi_stmt_2749: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2752_wire;
      req(0) <= phi_stmt_2749_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2749",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2749_ack_0,
          idata => idata,
          odata => conv797x_xlcssa_2749,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2749
    phi_stmt_2844: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2848_wire_constant & type_cast_2850_wire;
      req <= phi_stmt_2844_req_0 & phi_stmt_2844_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2844",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2844_ack_0,
          idata => idata,
          odata => k830x_x1_2844,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2844
    phi_stmt_2851: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2854_wire & type_cast_2856_wire;
      req <= phi_stmt_2851_req_0 & phi_stmt_2851_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2851",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2851_ack_0,
          idata => idata,
          odata => i834x_x2_2851,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2851
    phi_stmt_2857: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2861_wire_constant & type_cast_2863_wire;
      req <= phi_stmt_2857_req_0 & phi_stmt_2857_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2857",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2857_ack_0,
          idata => idata,
          odata => j884x_x1_2857,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2857
    phi_stmt_3262: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3266_wire_constant & type_cast_3268_wire;
      req <= phi_stmt_3262_req_0 & phi_stmt_3262_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3262",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3262_ack_0,
          idata => idata,
          odata => k830x_x0x_xph_3262,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3262
    phi_stmt_3269: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3272_wire & type_cast_3274_wire;
      req <= phi_stmt_3269_req_0 & phi_stmt_3269_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3269",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3269_ack_0,
          idata => idata,
          odata => i834x_x1x_xph_3269,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3269
    phi_stmt_3275: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3278_wire & type_cast_3280_wire;
      req <= phi_stmt_3275_req_0 & phi_stmt_3275_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3275",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3275_ack_0,
          idata => idata,
          odata => j884x_x0x_xph_3275,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3275
    phi_stmt_3284: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3287_wire;
      req(0) <= phi_stmt_3284_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3284",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3284_ack_0,
          idata => idata,
          odata => tmp1030x_xlcssa_3284,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3284
    phi_stmt_3288: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3291_wire;
      req(0) <= phi_stmt_3288_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3288",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3288_ack_0,
          idata => idata,
          odata => conv1015x_xlcssa_3288,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3288
    phi_stmt_3292: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3295_wire;
      req(0) <= phi_stmt_3292_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3292",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3292_ack_0,
          idata => idata,
          odata => tmp1014x_xlcssa_3292,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3292
    phi_stmt_3397: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3401_wire_constant & type_cast_3403_wire;
      req <= phi_stmt_3397_req_0 & phi_stmt_3397_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3397",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3397_ack_0,
          idata => idata,
          odata => k1050x_x1_3397,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3397
    phi_stmt_3404: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3407_wire & type_cast_3409_wire;
      req <= phi_stmt_3404_req_0 & phi_stmt_3404_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3404",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3404_ack_0,
          idata => idata,
          odata => i1058x_x2_3404,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3404
    phi_stmt_3410: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3413_wire & type_cast_3415_wire;
      req <= phi_stmt_3410_req_0 & phi_stmt_3410_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3410",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3410_ack_0,
          idata => idata,
          odata => j1108x_x1_3410,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3410
    phi_stmt_3801: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3804_wire & type_cast_3807_wire_constant;
      req <= phi_stmt_3801_req_0 & phi_stmt_3801_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3801",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3801_ack_0,
          idata => idata,
          odata => k1050x_x0x_xph_3801,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3801
    phi_stmt_3808: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3811_wire & type_cast_3813_wire;
      req <= phi_stmt_3808_req_0 & phi_stmt_3808_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3808",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3808_ack_0,
          idata => idata,
          odata => i1058x_x1x_xph_3808,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3808
    phi_stmt_3814: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3817_wire & type_cast_3819_wire;
      req <= phi_stmt_3814_req_0 & phi_stmt_3814_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3814",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3814_ack_0,
          idata => idata,
          odata => j1108x_x0x_xph_3814,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3814
    phi_stmt_3823: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3826_wire;
      req(0) <= phi_stmt_3823_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3823",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3823_ack_0,
          idata => idata,
          odata => tmp1252x_xlcssa_3823,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3823
    phi_stmt_3827: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_3830_wire;
      req(0) <= phi_stmt_3827_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3827",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3827_ack_0,
          idata => idata,
          odata => conv1238x_xlcssa_3827,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3827
    phi_stmt_3928: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3932_wire_constant & type_cast_3934_wire;
      req <= phi_stmt_3928_req_0 & phi_stmt_3928_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3928",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3928_ack_0,
          idata => idata,
          odata => k1272x_x1_3928,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3928
    phi_stmt_3935: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3938_wire & type_cast_3940_wire;
      req <= phi_stmt_3935_req_0 & phi_stmt_3935_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3935",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3935_ack_0,
          idata => idata,
          odata => i1276x_x2_3935,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3935
    phi_stmt_3941: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3945_wire_constant & type_cast_3947_wire;
      req <= phi_stmt_3941_req_0 & phi_stmt_3941_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3941",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3941_ack_0,
          idata => idata,
          odata => j1327x_x1_3941,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3941
    phi_stmt_4322: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4325_wire & type_cast_4328_wire_constant;
      req <= phi_stmt_4322_req_0 & phi_stmt_4322_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4322",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4322_ack_0,
          idata => idata,
          odata => k1272x_x0x_xph_4322,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4322
    phi_stmt_4329: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4332_wire & type_cast_4334_wire;
      req <= phi_stmt_4329_req_0 & phi_stmt_4329_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4329",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4329_ack_0,
          idata => idata,
          odata => i1276x_x1x_xph_4329,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4329
    phi_stmt_4335: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4338_wire & type_cast_4340_wire;
      req <= phi_stmt_4335_req_0 & phi_stmt_4335_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4335",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4335_ack_0,
          idata => idata,
          odata => j1327x_x0x_xph_4335,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4335
    phi_stmt_4344: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_4347_wire;
      req(0) <= phi_stmt_4344_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4344",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4344_ack_0,
          idata => idata,
          odata => tmp1471x_xlcssa_4344,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4344
    phi_stmt_4348: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_4351_wire;
      req(0) <= phi_stmt_4348_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4348",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4348_ack_0,
          idata => idata,
          odata => conv1456x_xlcssa_4348,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4348
    phi_stmt_4352: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_4355_wire;
      req(0) <= phi_stmt_4352_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4352",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4352_ack_0,
          idata => idata,
          odata => tmp1455x_xlcssa_4352,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4352
    phi_stmt_4463: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4467_wire_constant & type_cast_4469_wire;
      req <= phi_stmt_4463_req_0 & phi_stmt_4463_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4463",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4463_ack_0,
          idata => idata,
          odata => k1489x_x1_4463,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4463
    phi_stmt_4470: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4473_wire & type_cast_4475_wire;
      req <= phi_stmt_4470_req_0 & phi_stmt_4470_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4470",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4470_ack_0,
          idata => idata,
          odata => i1497x_x2_4470,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4470
    phi_stmt_4476: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4479_wire & type_cast_4481_wire;
      req <= phi_stmt_4476_req_0 & phi_stmt_4476_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4476",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4476_ack_0,
          idata => idata,
          odata => j1548x_x1_4476,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4476
    phi_stmt_4843: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4847_wire_constant & type_cast_4849_wire;
      req <= phi_stmt_4843_req_0 & phi_stmt_4843_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4843",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4843_ack_0,
          idata => idata,
          odata => k1489x_x0x_xph_4843,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4843
    phi_stmt_4850: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4853_wire & type_cast_4855_wire;
      req <= phi_stmt_4850_req_0 & phi_stmt_4850_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4850",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4850_ack_0,
          idata => idata,
          odata => i1497x_x1x_xph_4850,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4850
    phi_stmt_4856: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4859_wire & type_cast_4861_wire;
      req <= phi_stmt_4856_req_0 & phi_stmt_4856_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4856",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4856_ack_0,
          idata => idata,
          odata => j1548x_x0x_xph_4856,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4856
    phi_stmt_747: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_751_wire_constant & type_cast_753_wire;
      req <= phi_stmt_747_req_0 & phi_stmt_747_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_747",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_747_ack_0,
          idata => idata,
          odata => jx_x1_747,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_747
    phi_stmt_754: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_758_wire_constant & type_cast_760_wire;
      req <= phi_stmt_754_req_0 & phi_stmt_754_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_754",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_754_ack_0,
          idata => idata,
          odata => ix_x2_754,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_754
    phi_stmt_761: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_765_wire_constant & type_cast_767_wire;
      req <= phi_stmt_761_req_0 & phi_stmt_761_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_761",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_761_ack_0,
          idata => idata,
          odata => kx_x1_761,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_761
    -- flow-through select operator MUX_1118_inst
    jx_x2_1119 <= type_cast_1116_wire_constant when (cmp150_1103(0) /=  '0') else inc_1075;
    -- flow-through select operator MUX_1632_inst
    j230x_x2_1633 <= div181_1195 when (cmp364_1618(0) /=  '0') else inc355_1596;
    -- flow-through select operator MUX_2159_inst
    j446x_x2_2160 <= type_cast_2157_wire_constant when (cmp582_2144(0) /=  '0') else inc572_2116;
    -- flow-through select operator MUX_2686_inst
    j668x_x2_2687 <= div615_2240 when (cmp802_2672(0) /=  '0') else inc793_2650;
    -- flow-through select operator MUX_3219_inst
    j884x_x2_3220 <= type_cast_3217_wire_constant when (cmp1021_3204(0) /=  '0') else inc1011_3176;
    -- flow-through select operator MUX_3758_inst
    j1108x_x2_3759 <= div1055_3306 when (cmp1243_3744(0) /=  '0') else inc1234_3722;
    -- flow-through select operator MUX_4291_inst
    j1327x_x2_4292 <= type_cast_4289_wire_constant when (cmp1462_4276(0) /=  '0') else inc1452_4248;
    -- flow-through select operator MUX_4812_inst
    j1548x_x2_4813 <= div1494_4366 when (cmp1681_4798(0) /=  '0') else inc1672_4776;
    addr_of_1004_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1004_final_reg_req_0;
      addr_of_1004_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1004_final_reg_req_1;
      addr_of_1004_final_reg_ack_1<= rack(0);
      addr_of_1004_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1004_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1003_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx121_1005,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1029_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1029_final_reg_req_0;
      addr_of_1029_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1029_final_reg_req_1;
      addr_of_1029_final_reg_ack_1<= rack(0);
      addr_of_1029_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1029_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1028_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx126_1030,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1442_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1442_final_reg_req_0;
      addr_of_1442_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1442_final_reg_req_1;
      addr_of_1442_final_reg_ack_1<= rack(0);
      addr_of_1442_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1442_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1441_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx289_1443,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1525_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1525_final_reg_req_0;
      addr_of_1525_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1525_final_reg_req_1;
      addr_of_1525_final_reg_ack_1<= rack(0);
      addr_of_1525_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1525_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1524_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx332_1526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1550_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1550_final_reg_req_0;
      addr_of_1550_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1550_final_reg_req_1;
      addr_of_1550_final_reg_ack_1<= rack(0);
      addr_of_1550_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1550_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1549_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx337_1551,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1962_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1962_final_reg_req_0;
      addr_of_1962_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1962_final_reg_req_1;
      addr_of_1962_final_reg_ack_1<= rack(0);
      addr_of_1962_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1962_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1961_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx506_1963,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2045_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2045_final_reg_req_0;
      addr_of_2045_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2045_final_reg_req_1;
      addr_of_2045_final_reg_ack_1<= rack(0);
      addr_of_2045_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2045_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2044_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx549_2046,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2070_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2070_final_reg_req_0;
      addr_of_2070_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2070_final_reg_req_1;
      addr_of_2070_final_reg_ack_1<= rack(0);
      addr_of_2070_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2070_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2069_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx554_2071,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2496_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2496_final_reg_req_0;
      addr_of_2496_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2496_final_reg_req_1;
      addr_of_2496_final_reg_ack_1<= rack(0);
      addr_of_2496_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2496_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2495_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx727_2497,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2579_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2579_final_reg_req_0;
      addr_of_2579_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2579_final_reg_req_1;
      addr_of_2579_final_reg_ack_1<= rack(0);
      addr_of_2579_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2579_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2578_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx770_2580,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2604_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2604_final_reg_req_0;
      addr_of_2604_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2604_final_reg_req_1;
      addr_of_2604_final_reg_ack_1<= rack(0);
      addr_of_2604_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2604_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2603_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx775_2605,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3022_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3022_final_reg_req_0;
      addr_of_3022_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3022_final_reg_req_1;
      addr_of_3022_final_reg_ack_1<= rack(0);
      addr_of_3022_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3022_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3021_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx945_3023,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3105_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3105_final_reg_req_0;
      addr_of_3105_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3105_final_reg_req_1;
      addr_of_3105_final_reg_ack_1<= rack(0);
      addr_of_3105_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3105_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3104_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx988_3106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3130_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3130_final_reg_req_0;
      addr_of_3130_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3130_final_reg_req_1;
      addr_of_3130_final_reg_ack_1<= rack(0);
      addr_of_3130_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3130_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3129_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx993_3131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3568_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3568_final_reg_req_0;
      addr_of_3568_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3568_final_reg_req_1;
      addr_of_3568_final_reg_ack_1<= rack(0);
      addr_of_3568_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3568_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3567_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1168_3569,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3651_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3651_final_reg_req_0;
      addr_of_3651_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3651_final_reg_req_1;
      addr_of_3651_final_reg_ack_1<= rack(0);
      addr_of_3651_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3651_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3650_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1211_3652,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3676_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3676_final_reg_req_0;
      addr_of_3676_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3676_final_reg_req_1;
      addr_of_3676_final_reg_ack_1<= rack(0);
      addr_of_3676_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3676_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3675_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1216_3677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4094_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4094_final_reg_req_0;
      addr_of_4094_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4094_final_reg_req_1;
      addr_of_4094_final_reg_ack_1<= rack(0);
      addr_of_4094_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4094_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4093_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1386_4095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4177_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4177_final_reg_req_0;
      addr_of_4177_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4177_final_reg_req_1;
      addr_of_4177_final_reg_ack_1<= rack(0);
      addr_of_4177_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4177_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4176_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1429_4178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4202_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4202_final_reg_req_0;
      addr_of_4202_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4202_final_reg_req_1;
      addr_of_4202_final_reg_ack_1<= rack(0);
      addr_of_4202_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4202_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4201_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1434_4203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4622_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4622_final_reg_req_0;
      addr_of_4622_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4622_final_reg_req_1;
      addr_of_4622_final_reg_ack_1<= rack(0);
      addr_of_4622_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4622_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4621_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1606_4623,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4705_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4705_final_reg_req_0;
      addr_of_4705_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4705_final_reg_req_1;
      addr_of_4705_final_reg_ack_1<= rack(0);
      addr_of_4705_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4705_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4704_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1649_4706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4730_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4730_final_reg_req_0;
      addr_of_4730_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4730_final_reg_req_1;
      addr_of_4730_final_reg_ack_1<= rack(0);
      addr_of_4730_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4730_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4729_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1654_4731,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_921_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_921_final_reg_req_0;
      addr_of_921_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_921_final_reg_req_1;
      addr_of_921_final_reg_ack_1<= rack(0);
      addr_of_921_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_921_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_920_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_922,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1012_inst
    process(add117_984) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add117_984(31 downto 0);
      type_cast_1012_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1017_inst
    process(ASHR_i32_i32_1016_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1016_wire(31 downto 0);
      shr124_1018 <= tmp_var; -- 
    end process;
    type_cast_1022_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1022_inst_req_0;
      type_cast_1022_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1022_inst_req_1;
      type_cast_1022_inst_ack_1<= rack(0);
      type_cast_1022_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1022_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1021_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom125_1023,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1040_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1040_inst_req_0;
      type_cast_1040_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1040_inst_req_1;
      type_cast_1040_inst_ack_1<= rack(0);
      type_cast_1040_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1040_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1039_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv129_1041,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1050_inst
    process(add130_1047) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add130_1047(31 downto 0);
      type_cast_1050_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1052_inst
    process(conv21_677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv21_677(31 downto 0);
      type_cast_1052_wire <= tmp_var; -- 
    end process;
    type_cast_1079_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1079_inst_req_0;
      type_cast_1079_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1079_inst_req_1;
      type_cast_1079_inst_ack_1<= rack(0);
      type_cast_1079_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1079_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1078_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_1080,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1086_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1086_inst_req_0;
      type_cast_1086_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1086_inst_req_1;
      type_cast_1086_inst_ack_1<= rack(0);
      type_cast_1086_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1086_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp144_1083,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1087,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1106_inst_req_0;
      type_cast_1106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1106_inst_req_1;
      type_cast_1106_inst_ack_1<= rack(0);
      type_cast_1106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp150_1103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc155_1107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1123_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1123_inst_req_0;
      type_cast_1123_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1123_inst_req_1;
      type_cast_1123_inst_ack_1<= rack(0);
      type_cast_1123_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1123_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1122_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_1124,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1130_inst_req_0;
      type_cast_1130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1130_inst_req_1;
      type_cast_1130_inst_ack_1<= rack(0);
      type_cast_1130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp159_1127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv160_1131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1158_inst_req_0;
      type_cast_1158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1158_inst_req_1;
      type_cast_1158_inst_ack_1<= rack(0);
      type_cast_1158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1158_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1160_inst_req_0;
      type_cast_1160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1160_inst_req_1;
      type_cast_1160_inst_ack_1<= rack(0);
      type_cast_1160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1119,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1160_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1164_inst_req_0;
      type_cast_1164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1164_inst_req_1;
      type_cast_1164_inst_ack_1<= rack(0);
      type_cast_1164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_754,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1164_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1166_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1166_inst_req_0;
      type_cast_1166_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1166_inst_req_1;
      type_cast_1166_inst_ack_1<= rack(0);
      type_cast_1166_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1166_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc155x_xix_x2_1112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1166_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1170_inst_req_0;
      type_cast_1170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1170_inst_req_1;
      type_cast_1170_inst_ack_1<= rack(0);
      type_cast_1170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add138_1067,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1170_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1180_inst_req_0;
      type_cast_1180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1180_inst_req_1;
      type_cast_1180_inst_ack_1<= rack(0);
      type_cast_1180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv145_1087,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1180_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1184_inst_req_0;
      type_cast_1184_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1184_inst_req_1;
      type_cast_1184_inst_ack_1<= rack(0);
      type_cast_1184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp144_1083,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1184_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1188_inst_req_0;
      type_cast_1188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1188_inst_req_1;
      type_cast_1188_inst_ack_1<= rack(0);
      type_cast_1188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp144x_xlcssa_1181,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv180_1189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1210_inst_req_0;
      type_cast_1210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1210_inst_req_1;
      type_cast_1210_inst_ack_1<= rack(0);
      type_cast_1210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp191_1201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv216_1211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1214_inst_req_0;
      type_cast_1214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1214_inst_req_1;
      type_cast_1214_inst_ack_1<= rack(0);
      type_cast_1214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp203_1204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv224_1215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1218_inst_req_0;
      type_cast_1218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1218_inst_req_1;
      type_cast_1218_inst_ack_1<= rack(0);
      type_cast_1218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp207_1207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv226_1219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1227_inst_req_0;
      type_cast_1227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1227_inst_req_1;
      type_cast_1227_inst_ack_1<= rack(0);
      type_cast_1227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1227_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp187_1198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv238_1228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1231_inst_req_0;
      type_cast_1231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1231_inst_req_1;
      type_cast_1231_inst_ack_1<= rack(0);
      type_cast_1231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp203_1204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv275_1232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1241_inst
    process(sext1747_1238) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1747_1238(31 downto 0);
      type_cast_1241_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1246_inst
    process(ASHR_i32_i32_1245_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1245_wire(31 downto 0);
      conv281_1247 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1267_inst
    process(sext1707_1264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1707_1264(31 downto 0);
      type_cast_1267_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1272_inst
    process(ASHR_i32_i32_1271_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1271_wire(31 downto 0);
      conv305_1273 <= tmp_var; -- 
    end process;
    type_cast_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1279_inst_req_0;
      type_cast_1279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1279_inst_req_1;
      type_cast_1279_inst_ack_1<= rack(0);
      type_cast_1279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div181_1195,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1279_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1281_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1281_inst_req_0;
      type_cast_1281_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1281_inst_req_1;
      type_cast_1281_inst_ack_1<= rack(0);
      type_cast_1281_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1281_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j230x_x0x_xph_1669,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1281_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1288_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1288_inst_req_0;
      type_cast_1288_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1288_inst_req_1;
      type_cast_1288_inst_ack_1<= rack(0);
      type_cast_1288_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1288_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i184x_x1x_xph_1675,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1288_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1295_inst_req_0;
      type_cast_1295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1295_inst_req_1;
      type_cast_1295_inst_ack_1<= rack(0);
      type_cast_1295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k176x_x0x_xph_1681,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1295_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1300_inst_req_0;
      type_cast_1300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1300_inst_req_1;
      type_cast_1300_inst_ack_1<= rack(0);
      type_cast_1300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1300_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1299_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv236_1301,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1304_inst
    process(conv236_1301) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv236_1301(31 downto 0);
      type_cast_1304_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1306_inst
    process(conv238_1228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv238_1228(31 downto 0);
      type_cast_1306_wire <= tmp_var; -- 
    end process;
    type_cast_1321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1321_inst_req_0;
      type_cast_1321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1321_inst_req_1;
      type_cast_1321_inst_ack_1<= rack(0);
      type_cast_1321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp244_1318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv245_1322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1336_inst
    process(conv236_1301) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv236_1301(31 downto 0);
      type_cast_1336_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1338_inst
    process(add249_1333) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add249_1333(31 downto 0);
      type_cast_1338_wire <= tmp_var; -- 
    end process;
    type_cast_1351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1351_inst_req_0;
      type_cast_1351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1351_inst_req_1;
      type_cast_1351_inst_ack_1<= rack(0);
      type_cast_1351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1350_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv254_1352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1355_inst
    process(conv254_1352) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv254_1352(31 downto 0);
      type_cast_1355_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1357_inst
    process(conv238_1228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv238_1228(31 downto 0);
      type_cast_1357_wire <= tmp_var; -- 
    end process;
    type_cast_1372_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1372_inst_req_0;
      type_cast_1372_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1372_inst_req_1;
      type_cast_1372_inst_ack_1<= rack(0);
      type_cast_1372_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1372_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp262_1369,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv263_1373,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1381_inst
    process(conv254_1352) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv254_1352(31 downto 0);
      type_cast_1381_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1383_inst
    process(add266_1378) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add266_1378(31 downto 0);
      type_cast_1383_wire <= tmp_var; -- 
    end process;
    type_cast_1396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1396_inst_req_0;
      type_cast_1396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1396_inst_req_1;
      type_cast_1396_inst_ack_1<= rack(0);
      type_cast_1396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1395_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv273_1397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1401_inst_req_0;
      type_cast_1401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1401_inst_req_1;
      type_cast_1401_inst_ack_1<= rack(0);
      type_cast_1401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1400_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv277_1402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1425_inst
    process(add285_1422) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add285_1422(31 downto 0);
      type_cast_1425_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1430_inst
    process(ASHR_i32_i32_1429_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1429_wire(31 downto 0);
      shr287_1431 <= tmp_var; -- 
    end process;
    type_cast_1435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1435_inst_req_0;
      type_cast_1435_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1435_inst_req_1;
      type_cast_1435_inst_ack_1<= rack(0);
      type_cast_1435_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1435_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1434_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom288_1436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1454_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1454_inst_req_0;
      type_cast_1454_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1454_inst_req_1;
      type_cast_1454_inst_ack_1<= rack(0);
      type_cast_1454_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1454_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1453_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv294_1455,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1508_inst
    process(add312_1485) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add312_1485(31 downto 0);
      type_cast_1508_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1513_inst
    process(ASHR_i32_i32_1512_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1512_wire(31 downto 0);
      shr330_1514 <= tmp_var; -- 
    end process;
    type_cast_1518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1518_inst_req_0;
      type_cast_1518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1518_inst_req_1;
      type_cast_1518_inst_ack_1<= rack(0);
      type_cast_1518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1517_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom331_1519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1533_inst
    process(add328_1505) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add328_1505(31 downto 0);
      type_cast_1533_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1538_inst
    process(ASHR_i32_i32_1537_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1537_wire(31 downto 0);
      shr335_1539 <= tmp_var; -- 
    end process;
    type_cast_1543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1543_inst_req_0;
      type_cast_1543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1543_inst_req_1;
      type_cast_1543_inst_ack_1<= rack(0);
      type_cast_1543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1542_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom336_1544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1561_inst_req_0;
      type_cast_1561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1561_inst_req_1;
      type_cast_1561_inst_ack_1<= rack(0);
      type_cast_1561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1560_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv342_1562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1571_inst
    process(add343_1568) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add343_1568(31 downto 0);
      type_cast_1571_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1573_inst
    process(conv216_1211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv216_1211(31 downto 0);
      type_cast_1573_wire <= tmp_var; -- 
    end process;
    type_cast_1600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1600_inst_req_0;
      type_cast_1600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1600_inst_req_1;
      type_cast_1600_inst_ack_1<= rack(0);
      type_cast_1600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1599_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv357_1601,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1607_inst_req_0;
      type_cast_1607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1607_inst_req_1;
      type_cast_1607_inst_ack_1<= rack(0);
      type_cast_1607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp358_1604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv359_1608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1621_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1621_inst_req_0;
      type_cast_1621_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1621_inst_req_1;
      type_cast_1621_inst_ack_1<= rack(0);
      type_cast_1621_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1621_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp364_1618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc369_1622,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1637_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1637_inst_req_0;
      type_cast_1637_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1637_inst_req_1;
      type_cast_1637_inst_ack_1<= rack(0);
      type_cast_1637_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1637_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1636_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv372_1638,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1644_inst_req_0;
      type_cast_1644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1644_inst_req_1;
      type_cast_1644_inst_ack_1<= rack(0);
      type_cast_1644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp373_1641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv374_1645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1672_inst_req_0;
      type_cast_1672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1672_inst_req_1;
      type_cast_1672_inst_ack_1<= rack(0);
      type_cast_1672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1672_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j230x_x1_1276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1672_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1674_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1674_inst_req_0;
      type_cast_1674_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1674_inst_req_1;
      type_cast_1674_inst_ack_1<= rack(0);
      type_cast_1674_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1674_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j230x_x2_1633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1674_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1678_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1678_inst_req_0;
      type_cast_1678_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1678_inst_req_1;
      type_cast_1678_inst_ack_1<= rack(0);
      type_cast_1678_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1678_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc369x_xi184x_x2_1627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1678_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1680_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1680_inst_req_0;
      type_cast_1680_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1680_inst_req_1;
      type_cast_1680_inst_ack_1<= rack(0);
      type_cast_1680_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1680_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i184x_x2_1282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1680_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1684_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1684_inst_req_0;
      type_cast_1684_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1684_inst_req_1;
      type_cast_1684_inst_ack_1<= rack(0);
      type_cast_1684_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1684_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add351_1588,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1684_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1694_inst_req_0;
      type_cast_1694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1694_inst_req_1;
      type_cast_1694_inst_ack_1<= rack(0);
      type_cast_1694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp373_1641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1694_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1698_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1698_inst_req_0;
      type_cast_1698_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1698_inst_req_1;
      type_cast_1698_inst_ack_1<= rack(0);
      type_cast_1698_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1698_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv359_1608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1698_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1702_inst_req_0;
      type_cast_1702_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1702_inst_req_1;
      type_cast_1702_inst_ack_1<= rack(0);
      type_cast_1702_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1702_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp373x_xlcssa_1691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv398_1703,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1724_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1724_inst_req_0;
      type_cast_1724_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1724_inst_req_1;
      type_cast_1724_inst_ack_1<= rack(0);
      type_cast_1724_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1724_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp407_1715,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv432_1725,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1728_inst_req_0;
      type_cast_1728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1728_inst_req_1;
      type_cast_1728_inst_ack_1<= rack(0);
      type_cast_1728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp419_1718,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv440_1729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1732_inst_req_0;
      type_cast_1732_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1732_inst_req_1;
      type_cast_1732_inst_ack_1<= rack(0);
      type_cast_1732_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1732_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp423_1721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv442_1733,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1741_inst_req_0;
      type_cast_1741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1741_inst_req_1;
      type_cast_1741_inst_ack_1<= rack(0);
      type_cast_1741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp403_1712,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv454_1742,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1745_inst_req_0;
      type_cast_1745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1745_inst_req_1;
      type_cast_1745_inst_ack_1<= rack(0);
      type_cast_1745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp419_1718,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv492_1746,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1755_inst
    process(sext1748_1752) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1748_1752(31 downto 0);
      type_cast_1755_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1760_inst
    process(ASHR_i32_i32_1759_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1759_wire(31 downto 0);
      conv498_1761 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1781_inst
    process(sext1708_1778) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1708_1778(31 downto 0);
      type_cast_1781_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1786_inst
    process(ASHR_i32_i32_1785_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1785_wire(31 downto 0);
      conv522_1787 <= tmp_var; -- 
    end process;
    type_cast_1793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1793_inst_req_0;
      type_cast_1793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1793_inst_req_1;
      type_cast_1793_inst_ack_1<= rack(0);
      type_cast_1793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k392x_x0x_xph_2196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1793_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1800_inst_req_0;
      type_cast_1800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1800_inst_req_1;
      type_cast_1800_inst_ack_1<= rack(0);
      type_cast_1800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div399_1709,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1800_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1802_inst_req_0;
      type_cast_1802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1802_inst_req_1;
      type_cast_1802_inst_ack_1<= rack(0);
      type_cast_1802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i396x_x1x_xph_2203,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1802_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1809_inst_req_0;
      type_cast_1809_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1809_inst_req_1;
      type_cast_1809_inst_ack_1<= rack(0);
      type_cast_1809_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j446x_x0x_xph_2209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1809_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1814_inst_req_0;
      type_cast_1814_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1814_inst_req_1;
      type_cast_1814_inst_ack_1<= rack(0);
      type_cast_1814_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1814_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1813_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv452_1815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1818_inst
    process(conv452_1815) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv452_1815(31 downto 0);
      type_cast_1818_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1820_inst
    process(conv454_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv454_1742(31 downto 0);
      type_cast_1820_wire <= tmp_var; -- 
    end process;
    type_cast_1835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1835_inst_req_0;
      type_cast_1835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1835_inst_req_1;
      type_cast_1835_inst_ack_1<= rack(0);
      type_cast_1835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp460_1832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv461_1836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1850_inst
    process(conv452_1815) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv452_1815(31 downto 0);
      type_cast_1850_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1852_inst
    process(add465_1847) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add465_1847(31 downto 0);
      type_cast_1852_wire <= tmp_var; -- 
    end process;
    type_cast_1865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1865_inst_req_0;
      type_cast_1865_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1865_inst_req_1;
      type_cast_1865_inst_ack_1<= rack(0);
      type_cast_1865_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1864_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv470_1866,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1869_inst
    process(conv470_1866) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv470_1866(31 downto 0);
      type_cast_1869_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1871_inst
    process(conv454_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv454_1742(31 downto 0);
      type_cast_1871_wire <= tmp_var; -- 
    end process;
    type_cast_1886_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1886_inst_req_0;
      type_cast_1886_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1886_inst_req_1;
      type_cast_1886_inst_ack_1<= rack(0);
      type_cast_1886_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1886_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp478_1883,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv479_1887,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1901_inst
    process(conv470_1866) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv470_1866(31 downto 0);
      type_cast_1901_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1903_inst
    process(add483_1898) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add483_1898(31 downto 0);
      type_cast_1903_wire <= tmp_var; -- 
    end process;
    type_cast_1916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1916_inst_req_0;
      type_cast_1916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1916_inst_req_1;
      type_cast_1916_inst_ack_1<= rack(0);
      type_cast_1916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1915_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv490_1917,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1921_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1921_inst_req_0;
      type_cast_1921_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1921_inst_req_1;
      type_cast_1921_inst_ack_1<= rack(0);
      type_cast_1921_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1921_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1920_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv494_1922,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1945_inst
    process(add502_1942) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add502_1942(31 downto 0);
      type_cast_1945_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1950_inst
    process(ASHR_i32_i32_1949_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1949_wire(31 downto 0);
      shr504_1951 <= tmp_var; -- 
    end process;
    type_cast_1955_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1955_inst_req_0;
      type_cast_1955_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1955_inst_req_1;
      type_cast_1955_inst_ack_1<= rack(0);
      type_cast_1955_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1955_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1954_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom505_1956,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1974_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1974_inst_req_0;
      type_cast_1974_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1974_inst_req_1;
      type_cast_1974_inst_ack_1<= rack(0);
      type_cast_1974_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1974_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1973_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv511_1975,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2028_inst
    process(add529_2005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add529_2005(31 downto 0);
      type_cast_2028_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2033_inst
    process(ASHR_i32_i32_2032_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2032_wire(31 downto 0);
      shr547_2034 <= tmp_var; -- 
    end process;
    type_cast_2038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2038_inst_req_0;
      type_cast_2038_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2038_inst_req_1;
      type_cast_2038_inst_ack_1<= rack(0);
      type_cast_2038_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2037_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom548_2039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2053_inst
    process(add545_2025) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add545_2025(31 downto 0);
      type_cast_2053_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2058_inst
    process(ASHR_i32_i32_2057_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2057_wire(31 downto 0);
      shr552_2059 <= tmp_var; -- 
    end process;
    type_cast_2063_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2063_inst_req_0;
      type_cast_2063_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2063_inst_req_1;
      type_cast_2063_inst_ack_1<= rack(0);
      type_cast_2063_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2063_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2062_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom553_2064,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2081_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2081_inst_req_0;
      type_cast_2081_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2081_inst_req_1;
      type_cast_2081_inst_ack_1<= rack(0);
      type_cast_2081_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2081_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2080_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv559_2082,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2091_inst
    process(add560_2088) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add560_2088(31 downto 0);
      type_cast_2091_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2093_inst
    process(conv432_1725) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv432_1725(31 downto 0);
      type_cast_2093_wire <= tmp_var; -- 
    end process;
    type_cast_2120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2120_inst_req_0;
      type_cast_2120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2120_inst_req_1;
      type_cast_2120_inst_ack_1<= rack(0);
      type_cast_2120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2119_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv574_2121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2127_inst_req_0;
      type_cast_2127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2127_inst_req_1;
      type_cast_2127_inst_ack_1<= rack(0);
      type_cast_2127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp575_2124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv576_2128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2147_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2147_inst_req_0;
      type_cast_2147_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2147_inst_req_1;
      type_cast_2147_inst_ack_1<= rack(0);
      type_cast_2147_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2147_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp582_2144,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc587_2148,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2164_inst_req_0;
      type_cast_2164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2164_inst_req_1;
      type_cast_2164_inst_ack_1<= rack(0);
      type_cast_2164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2163_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv590_2165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2171_inst_req_0;
      type_cast_2171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2171_inst_req_1;
      type_cast_2171_inst_ack_1<= rack(0);
      type_cast_2171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2171_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp591_2168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv592_2172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2199_inst_req_0;
      type_cast_2199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2199_inst_req_1;
      type_cast_2199_inst_ack_1<= rack(0);
      type_cast_2199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add568_2108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2199_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2206_inst_req_0;
      type_cast_2206_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2206_inst_req_1;
      type_cast_2206_inst_ack_1<= rack(0);
      type_cast_2206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc587x_xi396x_x2_2153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2206_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2208_inst_req_0;
      type_cast_2208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2208_inst_req_1;
      type_cast_2208_inst_ack_1<= rack(0);
      type_cast_2208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i396x_x2_1797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2208_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2212_inst_req_0;
      type_cast_2212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2212_inst_req_1;
      type_cast_2212_inst_ack_1<= rack(0);
      type_cast_2212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j446x_x2_2160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2212_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2214_inst_req_0;
      type_cast_2214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2214_inst_req_1;
      type_cast_2214_inst_ack_1<= rack(0);
      type_cast_2214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j446x_x1_1803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2214_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2221_inst_req_0;
      type_cast_2221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2221_inst_req_1;
      type_cast_2221_inst_ack_1<= rack(0);
      type_cast_2221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp591_2168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2221_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2225_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2225_inst_req_0;
      type_cast_2225_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2225_inst_req_1;
      type_cast_2225_inst_ack_1<= rack(0);
      type_cast_2225_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2225_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv576_2128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2225_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2229_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2229_inst_req_0;
      type_cast_2229_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2229_inst_req_1;
      type_cast_2229_inst_ack_1<= rack(0);
      type_cast_2229_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2229_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp575_2124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2229_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2233_inst_req_0;
      type_cast_2233_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2233_inst_req_1;
      type_cast_2233_inst_ack_1<= rack(0);
      type_cast_2233_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp575x_xlcssa_2226,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv614_2234,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2243_inst_req_0;
      type_cast_2243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2243_inst_req_1;
      type_cast_2243_inst_ack_1<= rack(0);
      type_cast_2243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp591x_xlcssa_2218,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv620_2244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2265_inst_req_0;
      type_cast_2265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2265_inst_req_1;
      type_cast_2265_inst_ack_1<= rack(0);
      type_cast_2265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp629_2256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv654_2266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2269_inst_req_0;
      type_cast_2269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2269_inst_req_1;
      type_cast_2269_inst_ack_1<= rack(0);
      type_cast_2269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp641_2259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv662_2270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2273_inst_req_0;
      type_cast_2273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2273_inst_req_1;
      type_cast_2273_inst_ack_1<= rack(0);
      type_cast_2273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp645_2262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv664_2274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2282_inst_req_0;
      type_cast_2282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2282_inst_req_1;
      type_cast_2282_inst_ack_1<= rack(0);
      type_cast_2282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp625_2253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv676_2283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2286_inst_req_0;
      type_cast_2286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2286_inst_req_1;
      type_cast_2286_inst_ack_1<= rack(0);
      type_cast_2286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp641_2259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv713_2287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2296_inst
    process(sext1749_2293) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1749_2293(31 downto 0);
      type_cast_2296_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2301_inst
    process(ASHR_i32_i32_2300_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2300_wire(31 downto 0);
      conv719_2302 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2322_inst
    process(sext1709_2319) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1709_2319(31 downto 0);
      type_cast_2322_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2327_inst
    process(ASHR_i32_i32_2326_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2326_wire(31 downto 0);
      conv743_2328 <= tmp_var; -- 
    end process;
    type_cast_2337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2337_inst_req_0;
      type_cast_2337_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2337_inst_req_1;
      type_cast_2337_inst_ack_1<= rack(0);
      type_cast_2337_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2337_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k610x_x0x_xph_2723,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2337_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2341_inst_req_0;
      type_cast_2341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2341_inst_req_1;
      type_cast_2341_inst_ack_1<= rack(0);
      type_cast_2341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div621_2250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2341_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2343_inst_req_0;
      type_cast_2343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2343_inst_req_1;
      type_cast_2343_inst_ack_1<= rack(0);
      type_cast_2343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i618x_x1x_xph_2730,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2343_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2347_inst_req_0;
      type_cast_2347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2347_inst_req_1;
      type_cast_2347_inst_ack_1<= rack(0);
      type_cast_2347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div615_2240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2347_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2349_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2349_inst_req_0;
      type_cast_2349_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2349_inst_req_1;
      type_cast_2349_inst_ack_1<= rack(0);
      type_cast_2349_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2349_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j668x_x0x_xph_2736,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2349_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2354_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2354_inst_req_0;
      type_cast_2354_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2354_inst_req_1;
      type_cast_2354_inst_ack_1<= rack(0);
      type_cast_2354_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2354_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2353_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv674_2355,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2358_inst
    process(conv674_2355) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv674_2355(31 downto 0);
      type_cast_2358_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2360_inst
    process(conv676_2283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv676_2283(31 downto 0);
      type_cast_2360_wire <= tmp_var; -- 
    end process;
    type_cast_2375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2375_inst_req_0;
      type_cast_2375_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2375_inst_req_1;
      type_cast_2375_inst_ack_1<= rack(0);
      type_cast_2375_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2375_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp682_2372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv683_2376,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2390_inst
    process(conv674_2355) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv674_2355(31 downto 0);
      type_cast_2390_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2392_inst
    process(add687_2387) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add687_2387(31 downto 0);
      type_cast_2392_wire <= tmp_var; -- 
    end process;
    type_cast_2405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2405_inst_req_0;
      type_cast_2405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2405_inst_req_1;
      type_cast_2405_inst_ack_1<= rack(0);
      type_cast_2405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2404_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv692_2406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2409_inst
    process(conv692_2406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv692_2406(31 downto 0);
      type_cast_2409_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2411_inst
    process(conv676_2283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv676_2283(31 downto 0);
      type_cast_2411_wire <= tmp_var; -- 
    end process;
    type_cast_2426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2426_inst_req_0;
      type_cast_2426_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2426_inst_req_1;
      type_cast_2426_inst_ack_1<= rack(0);
      type_cast_2426_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2426_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp700_2423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv701_2427,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2435_inst
    process(conv692_2406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv692_2406(31 downto 0);
      type_cast_2435_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2437_inst
    process(add704_2432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add704_2432(31 downto 0);
      type_cast_2437_wire <= tmp_var; -- 
    end process;
    type_cast_2450_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2450_inst_req_0;
      type_cast_2450_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2450_inst_req_1;
      type_cast_2450_inst_ack_1<= rack(0);
      type_cast_2450_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2450_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2449_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv711_2451,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2455_inst_req_0;
      type_cast_2455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2455_inst_req_1;
      type_cast_2455_inst_ack_1<= rack(0);
      type_cast_2455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2454_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv715_2456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2479_inst
    process(add723_2476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add723_2476(31 downto 0);
      type_cast_2479_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2484_inst
    process(ASHR_i32_i32_2483_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2483_wire(31 downto 0);
      shr725_2485 <= tmp_var; -- 
    end process;
    type_cast_2489_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2489_inst_req_0;
      type_cast_2489_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2489_inst_req_1;
      type_cast_2489_inst_ack_1<= rack(0);
      type_cast_2489_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2489_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2488_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom726_2490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2508_inst_req_0;
      type_cast_2508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2508_inst_req_1;
      type_cast_2508_inst_ack_1<= rack(0);
      type_cast_2508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2507_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv732_2509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2562_inst
    process(add750_2539) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add750_2539(31 downto 0);
      type_cast_2562_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2567_inst
    process(ASHR_i32_i32_2566_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2566_wire(31 downto 0);
      shr768_2568 <= tmp_var; -- 
    end process;
    type_cast_2572_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2572_inst_req_0;
      type_cast_2572_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2572_inst_req_1;
      type_cast_2572_inst_ack_1<= rack(0);
      type_cast_2572_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2572_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2571_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom769_2573,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2587_inst
    process(add766_2559) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add766_2559(31 downto 0);
      type_cast_2587_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2592_inst
    process(ASHR_i32_i32_2591_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2591_wire(31 downto 0);
      shr773_2593 <= tmp_var; -- 
    end process;
    type_cast_2597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2597_inst_req_0;
      type_cast_2597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2597_inst_req_1;
      type_cast_2597_inst_ack_1<= rack(0);
      type_cast_2597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2596_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom774_2598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2615_inst_req_0;
      type_cast_2615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2615_inst_req_1;
      type_cast_2615_inst_ack_1<= rack(0);
      type_cast_2615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2614_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv780_2616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2625_inst
    process(add781_2622) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add781_2622(31 downto 0);
      type_cast_2625_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2627_inst
    process(conv654_2266) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv654_2266(31 downto 0);
      type_cast_2627_wire <= tmp_var; -- 
    end process;
    type_cast_2654_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2654_inst_req_0;
      type_cast_2654_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2654_inst_req_1;
      type_cast_2654_inst_ack_1<= rack(0);
      type_cast_2654_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2654_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2653_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv795_2655,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2661_inst_req_0;
      type_cast_2661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2661_inst_req_1;
      type_cast_2661_inst_ack_1<= rack(0);
      type_cast_2661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp796_2658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv797_2662,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2675_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2675_inst_req_0;
      type_cast_2675_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2675_inst_req_1;
      type_cast_2675_inst_ack_1<= rack(0);
      type_cast_2675_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2675_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp802_2672,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc807_2676,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2691_inst_req_0;
      type_cast_2691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2691_inst_req_1;
      type_cast_2691_inst_ack_1<= rack(0);
      type_cast_2691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2690_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv810_2692,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2698_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2698_inst_req_0;
      type_cast_2698_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2698_inst_req_1;
      type_cast_2698_inst_ack_1<= rack(0);
      type_cast_2698_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2698_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp811_2695,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv812_2699,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2726_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2726_inst_req_0;
      type_cast_2726_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2726_inst_req_1;
      type_cast_2726_inst_ack_1<= rack(0);
      type_cast_2726_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2726_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add789_2642,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2726_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2733_inst_req_0;
      type_cast_2733_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2733_inst_req_1;
      type_cast_2733_inst_ack_1<= rack(0);
      type_cast_2733_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2733_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i618x_x2_2338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2733_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2735_inst_req_0;
      type_cast_2735_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2735_inst_req_1;
      type_cast_2735_inst_ack_1<= rack(0);
      type_cast_2735_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2735_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc807x_xi618x_x2_2681,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2735_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2739_inst_req_0;
      type_cast_2739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2739_inst_req_1;
      type_cast_2739_inst_ack_1<= rack(0);
      type_cast_2739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j668x_x1_2344,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2739_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2741_inst_req_0;
      type_cast_2741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2741_inst_req_1;
      type_cast_2741_inst_ack_1<= rack(0);
      type_cast_2741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j668x_x2_2687,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2741_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2748_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2748_inst_req_0;
      type_cast_2748_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2748_inst_req_1;
      type_cast_2748_inst_ack_1<= rack(0);
      type_cast_2748_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2748_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp811_2695,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2748_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2752_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2752_inst_req_0;
      type_cast_2752_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2752_inst_req_1;
      type_cast_2752_inst_ack_1<= rack(0);
      type_cast_2752_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2752_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv797_2662,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2752_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2756_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2756_inst_req_0;
      type_cast_2756_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2756_inst_req_1;
      type_cast_2756_inst_ack_1<= rack(0);
      type_cast_2756_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2756_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp811x_xlcssa_2745,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv836_2757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2778_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2778_inst_req_0;
      type_cast_2778_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2778_inst_req_1;
      type_cast_2778_inst_ack_1<= rack(0);
      type_cast_2778_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2778_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp845_2769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv870_2779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2782_inst_req_0;
      type_cast_2782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2782_inst_req_1;
      type_cast_2782_inst_ack_1<= rack(0);
      type_cast_2782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp857_2772,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv878_2783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2786_inst_req_0;
      type_cast_2786_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2786_inst_req_1;
      type_cast_2786_inst_ack_1<= rack(0);
      type_cast_2786_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2786_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp861_2775,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv880_2787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2795_inst_req_0;
      type_cast_2795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2795_inst_req_1;
      type_cast_2795_inst_ack_1<= rack(0);
      type_cast_2795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp841_2766,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv892_2796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2799_inst_req_0;
      type_cast_2799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2799_inst_req_1;
      type_cast_2799_inst_ack_1<= rack(0);
      type_cast_2799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp857_2772,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv931_2800,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2809_inst
    process(sext1750_2806) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1750_2806(31 downto 0);
      type_cast_2809_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2814_inst
    process(ASHR_i32_i32_2813_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2813_wire(31 downto 0);
      conv937_2815 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2835_inst
    process(sext1710_2832) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1710_2832(31 downto 0);
      type_cast_2835_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2840_inst
    process(ASHR_i32_i32_2839_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2839_wire(31 downto 0);
      conv961_2841 <= tmp_var; -- 
    end process;
    type_cast_2850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2850_inst_req_0;
      type_cast_2850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2850_inst_req_1;
      type_cast_2850_inst_ack_1<= rack(0);
      type_cast_2850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k830x_x0x_xph_3262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2850_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2854_inst_req_0;
      type_cast_2854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2854_inst_req_1;
      type_cast_2854_inst_ack_1<= rack(0);
      type_cast_2854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div837_2763,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2854_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2856_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2856_inst_req_0;
      type_cast_2856_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2856_inst_req_1;
      type_cast_2856_inst_ack_1<= rack(0);
      type_cast_2856_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2856_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i834x_x1x_xph_3269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2856_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2863_inst_req_0;
      type_cast_2863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2863_inst_req_1;
      type_cast_2863_inst_ack_1<= rack(0);
      type_cast_2863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j884x_x0x_xph_3275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2863_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2868_inst_req_0;
      type_cast_2868_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2868_inst_req_1;
      type_cast_2868_inst_ack_1<= rack(0);
      type_cast_2868_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2868_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2867_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv890_2869,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2872_inst
    process(conv890_2869) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv890_2869(31 downto 0);
      type_cast_2872_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2874_inst
    process(conv892_2796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv892_2796(31 downto 0);
      type_cast_2874_wire <= tmp_var; -- 
    end process;
    type_cast_2889_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2889_inst_req_0;
      type_cast_2889_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2889_inst_req_1;
      type_cast_2889_inst_ack_1<= rack(0);
      type_cast_2889_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2889_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp898_2886,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv899_2890,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2910_inst
    process(conv890_2869) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv890_2869(31 downto 0);
      type_cast_2910_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2912_inst
    process(add904_2907) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add904_2907(31 downto 0);
      type_cast_2912_wire <= tmp_var; -- 
    end process;
    type_cast_2925_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2925_inst_req_0;
      type_cast_2925_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2925_inst_req_1;
      type_cast_2925_inst_ack_1<= rack(0);
      type_cast_2925_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2925_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2924_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv909_2926,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2929_inst
    process(conv909_2926) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv909_2926(31 downto 0);
      type_cast_2929_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2931_inst
    process(conv892_2796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv892_2796(31 downto 0);
      type_cast_2931_wire <= tmp_var; -- 
    end process;
    type_cast_2946_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2946_inst_req_0;
      type_cast_2946_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2946_inst_req_1;
      type_cast_2946_inst_ack_1<= rack(0);
      type_cast_2946_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2946_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp917_2943,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv918_2947,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2961_inst
    process(conv909_2926) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv909_2926(31 downto 0);
      type_cast_2961_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2963_inst
    process(add922_2958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add922_2958(31 downto 0);
      type_cast_2963_wire <= tmp_var; -- 
    end process;
    type_cast_2976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2976_inst_req_0;
      type_cast_2976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2976_inst_req_1;
      type_cast_2976_inst_ack_1<= rack(0);
      type_cast_2976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2975_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv929_2977,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2981_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2981_inst_req_0;
      type_cast_2981_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2981_inst_req_1;
      type_cast_2981_inst_ack_1<= rack(0);
      type_cast_2981_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2981_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2980_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv933_2982,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3005_inst
    process(add941_3002) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add941_3002(31 downto 0);
      type_cast_3005_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3010_inst
    process(ASHR_i32_i32_3009_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3009_wire(31 downto 0);
      shr943_3011 <= tmp_var; -- 
    end process;
    type_cast_3015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3015_inst_req_0;
      type_cast_3015_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3015_inst_req_1;
      type_cast_3015_inst_ack_1<= rack(0);
      type_cast_3015_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3015_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3014_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom944_3016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3034_inst_req_0;
      type_cast_3034_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3034_inst_req_1;
      type_cast_3034_inst_ack_1<= rack(0);
      type_cast_3034_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3034_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3033_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv950_3035,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3088_inst
    process(add968_3065) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add968_3065(31 downto 0);
      type_cast_3088_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3093_inst
    process(ASHR_i32_i32_3092_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3092_wire(31 downto 0);
      shr986_3094 <= tmp_var; -- 
    end process;
    type_cast_3098_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3098_inst_req_0;
      type_cast_3098_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3098_inst_req_1;
      type_cast_3098_inst_ack_1<= rack(0);
      type_cast_3098_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3098_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3097_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom987_3099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3113_inst
    process(add984_3085) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add984_3085(31 downto 0);
      type_cast_3113_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3118_inst
    process(ASHR_i32_i32_3117_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3117_wire(31 downto 0);
      shr991_3119 <= tmp_var; -- 
    end process;
    type_cast_3123_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3123_inst_req_0;
      type_cast_3123_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3123_inst_req_1;
      type_cast_3123_inst_ack_1<= rack(0);
      type_cast_3123_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3123_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3122_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom992_3124,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3141_inst_req_0;
      type_cast_3141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3141_inst_req_1;
      type_cast_3141_inst_ack_1<= rack(0);
      type_cast_3141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3140_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv998_3142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3151_inst
    process(add999_3148) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add999_3148(31 downto 0);
      type_cast_3151_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3153_inst
    process(conv870_2779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv870_2779(31 downto 0);
      type_cast_3153_wire <= tmp_var; -- 
    end process;
    type_cast_3180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3180_inst_req_0;
      type_cast_3180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3180_inst_req_1;
      type_cast_3180_inst_ack_1<= rack(0);
      type_cast_3180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3179_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1013_3181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3187_inst_req_0;
      type_cast_3187_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3187_inst_req_1;
      type_cast_3187_inst_ack_1<= rack(0);
      type_cast_3187_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1014_3184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1015_3188,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3207_inst_req_0;
      type_cast_3207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3207_inst_req_1;
      type_cast_3207_inst_ack_1<= rack(0);
      type_cast_3207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1021_3204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1026_3208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3224_inst_req_0;
      type_cast_3224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3224_inst_req_1;
      type_cast_3224_inst_ack_1<= rack(0);
      type_cast_3224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3223_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1029_3225,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3231_inst_req_0;
      type_cast_3231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3231_inst_req_1;
      type_cast_3231_inst_ack_1<= rack(0);
      type_cast_3231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1030_3228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1031_3232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3268_inst_req_0;
      type_cast_3268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3268_inst_req_1;
      type_cast_3268_inst_ack_1<= rack(0);
      type_cast_3268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1007_3168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3268_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3272_inst_req_0;
      type_cast_3272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3272_inst_req_1;
      type_cast_3272_inst_ack_1<= rack(0);
      type_cast_3272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i834x_x2_2851,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3272_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3274_inst_req_0;
      type_cast_3274_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3274_inst_req_1;
      type_cast_3274_inst_ack_1<= rack(0);
      type_cast_3274_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3274_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1026x_xi834x_x2_3213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3274_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3278_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3278_inst_req_0;
      type_cast_3278_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3278_inst_req_1;
      type_cast_3278_inst_ack_1<= rack(0);
      type_cast_3278_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3278_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j884x_x2_3220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3278_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3280_inst_req_0;
      type_cast_3280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3280_inst_req_1;
      type_cast_3280_inst_ack_1<= rack(0);
      type_cast_3280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j884x_x1_2857,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3280_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3287_inst_req_0;
      type_cast_3287_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3287_inst_req_1;
      type_cast_3287_inst_ack_1<= rack(0);
      type_cast_3287_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3287_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1030_3228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3287_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3291_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3291_inst_req_0;
      type_cast_3291_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3291_inst_req_1;
      type_cast_3291_inst_ack_1<= rack(0);
      type_cast_3291_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3291_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv1015_3188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3291_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3295_inst_req_0;
      type_cast_3295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3295_inst_req_1;
      type_cast_3295_inst_ack_1<= rack(0);
      type_cast_3295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1014_3184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3295_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3299_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3299_inst_req_0;
      type_cast_3299_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3299_inst_req_1;
      type_cast_3299_inst_ack_1<= rack(0);
      type_cast_3299_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3299_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1014x_xlcssa_3292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1054_3300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3309_inst_req_0;
      type_cast_3309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3309_inst_req_1;
      type_cast_3309_inst_ack_1<= rack(0);
      type_cast_3309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1030x_xlcssa_3284,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1060_3310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3331_inst_req_0;
      type_cast_3331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3331_inst_req_1;
      type_cast_3331_inst_ack_1<= rack(0);
      type_cast_3331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1069_3322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1094_3332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3335_inst_req_0;
      type_cast_3335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3335_inst_req_1;
      type_cast_3335_inst_ack_1<= rack(0);
      type_cast_3335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3335_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1081_3325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1102_3336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3339_inst_req_0;
      type_cast_3339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3339_inst_req_1;
      type_cast_3339_inst_ack_1<= rack(0);
      type_cast_3339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1085_3328,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1104_3340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3348_inst_req_0;
      type_cast_3348_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3348_inst_req_1;
      type_cast_3348_inst_ack_1<= rack(0);
      type_cast_3348_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1065_3319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1116_3349,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3352_inst_req_0;
      type_cast_3352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3352_inst_req_1;
      type_cast_3352_inst_ack_1<= rack(0);
      type_cast_3352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1081_3325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1154_3353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3362_inst
    process(sext1751_3359) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1751_3359(31 downto 0);
      type_cast_3362_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3367_inst
    process(ASHR_i32_i32_3366_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3366_wire(31 downto 0);
      conv1160_3368 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3388_inst
    process(sext1711_3385) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1711_3385(31 downto 0);
      type_cast_3388_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3393_inst
    process(ASHR_i32_i32_3392_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3392_wire(31 downto 0);
      conv1184_3394 <= tmp_var; -- 
    end process;
    type_cast_3403_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3403_inst_req_0;
      type_cast_3403_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3403_inst_req_1;
      type_cast_3403_inst_ack_1<= rack(0);
      type_cast_3403_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3403_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1050x_x0x_xph_3801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3403_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3407_inst_req_0;
      type_cast_3407_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3407_inst_req_1;
      type_cast_3407_inst_ack_1<= rack(0);
      type_cast_3407_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3407_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1058x_x1x_xph_3808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3407_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3409_inst_req_0;
      type_cast_3409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3409_inst_req_1;
      type_cast_3409_inst_ack_1<= rack(0);
      type_cast_3409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1061_3316,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3409_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3413_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3413_inst_req_0;
      type_cast_3413_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3413_inst_req_1;
      type_cast_3413_inst_ack_1<= rack(0);
      type_cast_3413_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3413_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1055_3306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3413_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3415_inst_req_0;
      type_cast_3415_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3415_inst_req_1;
      type_cast_3415_inst_ack_1<= rack(0);
      type_cast_3415_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3415_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1108x_x0x_xph_3814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3415_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3420_inst_req_0;
      type_cast_3420_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3420_inst_req_1;
      type_cast_3420_inst_ack_1<= rack(0);
      type_cast_3420_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3420_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3419_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1114_3421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3424_inst
    process(conv1114_3421) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1114_3421(31 downto 0);
      type_cast_3424_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3426_inst
    process(conv1116_3349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1116_3349(31 downto 0);
      type_cast_3426_wire <= tmp_var; -- 
    end process;
    type_cast_3441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3441_inst_req_0;
      type_cast_3441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3441_inst_req_1;
      type_cast_3441_inst_ack_1<= rack(0);
      type_cast_3441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1122_3438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1123_3442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3462_inst
    process(conv1114_3421) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1114_3421(31 downto 0);
      type_cast_3462_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3464_inst
    process(add1128_3459) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1128_3459(31 downto 0);
      type_cast_3464_wire <= tmp_var; -- 
    end process;
    type_cast_3477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3477_inst_req_0;
      type_cast_3477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3477_inst_req_1;
      type_cast_3477_inst_ack_1<= rack(0);
      type_cast_3477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3476_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1133_3478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3481_inst
    process(conv1133_3478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1133_3478(31 downto 0);
      type_cast_3481_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3483_inst
    process(conv1116_3349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1116_3349(31 downto 0);
      type_cast_3483_wire <= tmp_var; -- 
    end process;
    type_cast_3498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3498_inst_req_0;
      type_cast_3498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3498_inst_req_1;
      type_cast_3498_inst_ack_1<= rack(0);
      type_cast_3498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1141_3495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1142_3499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3507_inst
    process(conv1133_3478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1133_3478(31 downto 0);
      type_cast_3507_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3509_inst
    process(add1145_3504) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1145_3504(31 downto 0);
      type_cast_3509_wire <= tmp_var; -- 
    end process;
    type_cast_3522_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3522_inst_req_0;
      type_cast_3522_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3522_inst_req_1;
      type_cast_3522_inst_ack_1<= rack(0);
      type_cast_3522_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3522_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3521_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1152_3523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3527_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3527_inst_req_0;
      type_cast_3527_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3527_inst_req_1;
      type_cast_3527_inst_ack_1<= rack(0);
      type_cast_3527_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3527_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3526_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1156_3528,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3551_inst
    process(add1164_3548) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1164_3548(31 downto 0);
      type_cast_3551_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3556_inst
    process(ASHR_i32_i32_3555_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3555_wire(31 downto 0);
      shr1166_3557 <= tmp_var; -- 
    end process;
    type_cast_3561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3561_inst_req_0;
      type_cast_3561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3561_inst_req_1;
      type_cast_3561_inst_ack_1<= rack(0);
      type_cast_3561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3560_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1167_3562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3580_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3580_inst_req_0;
      type_cast_3580_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3580_inst_req_1;
      type_cast_3580_inst_ack_1<= rack(0);
      type_cast_3580_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3580_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3579_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1173_3581,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3634_inst
    process(add1191_3611) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1191_3611(31 downto 0);
      type_cast_3634_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3639_inst
    process(ASHR_i32_i32_3638_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3638_wire(31 downto 0);
      shr1209_3640 <= tmp_var; -- 
    end process;
    type_cast_3644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3644_inst_req_0;
      type_cast_3644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3644_inst_req_1;
      type_cast_3644_inst_ack_1<= rack(0);
      type_cast_3644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3643_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1210_3645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3659_inst
    process(add1207_3631) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1207_3631(31 downto 0);
      type_cast_3659_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3664_inst
    process(ASHR_i32_i32_3663_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3663_wire(31 downto 0);
      shr1214_3665 <= tmp_var; -- 
    end process;
    type_cast_3669_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3669_inst_req_0;
      type_cast_3669_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3669_inst_req_1;
      type_cast_3669_inst_ack_1<= rack(0);
      type_cast_3669_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3669_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3668_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1215_3670,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3687_inst_req_0;
      type_cast_3687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3687_inst_req_1;
      type_cast_3687_inst_ack_1<= rack(0);
      type_cast_3687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3686_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1221_3688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3697_inst
    process(add1222_3694) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1222_3694(31 downto 0);
      type_cast_3697_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3699_inst
    process(conv1094_3332) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1094_3332(31 downto 0);
      type_cast_3699_wire <= tmp_var; -- 
    end process;
    type_cast_3726_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3726_inst_req_0;
      type_cast_3726_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3726_inst_req_1;
      type_cast_3726_inst_ack_1<= rack(0);
      type_cast_3726_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3726_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3725_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1236_3727,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3733_inst_req_0;
      type_cast_3733_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3733_inst_req_1;
      type_cast_3733_inst_ack_1<= rack(0);
      type_cast_3733_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3733_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1237_3730,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1238_3734,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3747_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3747_inst_req_0;
      type_cast_3747_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3747_inst_req_1;
      type_cast_3747_inst_ack_1<= rack(0);
      type_cast_3747_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3747_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1243_3744,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1248_3748,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3763_inst_req_0;
      type_cast_3763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3763_inst_req_1;
      type_cast_3763_inst_ack_1<= rack(0);
      type_cast_3763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3762_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1251_3764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3770_inst_req_0;
      type_cast_3770_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3770_inst_req_1;
      type_cast_3770_inst_ack_1<= rack(0);
      type_cast_3770_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3770_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1252_3767,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1253_3771,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3804_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3804_inst_req_0;
      type_cast_3804_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3804_inst_req_1;
      type_cast_3804_inst_ack_1<= rack(0);
      type_cast_3804_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3804_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1230_3714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3804_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3811_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3811_inst_req_0;
      type_cast_3811_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3811_inst_req_1;
      type_cast_3811_inst_ack_1<= rack(0);
      type_cast_3811_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3811_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1058x_x2_3404,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3811_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3813_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3813_inst_req_0;
      type_cast_3813_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3813_inst_req_1;
      type_cast_3813_inst_ack_1<= rack(0);
      type_cast_3813_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3813_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1248x_xi1058x_x2_3753,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3813_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3817_inst_req_0;
      type_cast_3817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3817_inst_req_1;
      type_cast_3817_inst_ack_1<= rack(0);
      type_cast_3817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1108x_x1_3410,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3817_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3819_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3819_inst_req_0;
      type_cast_3819_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3819_inst_req_1;
      type_cast_3819_inst_ack_1<= rack(0);
      type_cast_3819_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3819_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1108x_x2_3759,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3819_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3826_inst_req_0;
      type_cast_3826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3826_inst_req_1;
      type_cast_3826_inst_ack_1<= rack(0);
      type_cast_3826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1252_3767,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3826_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3830_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3830_inst_req_0;
      type_cast_3830_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3830_inst_req_1;
      type_cast_3830_inst_ack_1<= rack(0);
      type_cast_3830_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3830_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv1238_3734,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3830_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3834_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3834_inst_req_0;
      type_cast_3834_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3834_inst_req_1;
      type_cast_3834_inst_ack_1<= rack(0);
      type_cast_3834_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3834_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1252x_xlcssa_3823,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1278_3835,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3862_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3862_inst_req_0;
      type_cast_3862_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3862_inst_req_1;
      type_cast_3862_inst_ack_1<= rack(0);
      type_cast_3862_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3862_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1288_3853,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1313_3863,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3866_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3866_inst_req_0;
      type_cast_3866_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3866_inst_req_1;
      type_cast_3866_inst_ack_1<= rack(0);
      type_cast_3866_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3866_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1300_3856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1321_3867,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3870_inst_req_0;
      type_cast_3870_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3870_inst_req_1;
      type_cast_3870_inst_ack_1<= rack(0);
      type_cast_3870_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1304_3859,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1323_3871,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3879_inst_req_0;
      type_cast_3879_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3879_inst_req_1;
      type_cast_3879_inst_ack_1<= rack(0);
      type_cast_3879_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3879_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1284_3850,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1335_3880,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3883_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3883_inst_req_0;
      type_cast_3883_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3883_inst_req_1;
      type_cast_3883_inst_ack_1<= rack(0);
      type_cast_3883_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3883_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1300_3856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1372_3884,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3893_inst
    process(sext1752_3890) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1752_3890(31 downto 0);
      type_cast_3893_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3898_inst
    process(ASHR_i32_i32_3897_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3897_wire(31 downto 0);
      conv1378_3899 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3919_inst
    process(sext1712_3916) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1712_3916(31 downto 0);
      type_cast_3919_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3924_inst
    process(ASHR_i32_i32_3923_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3923_wire(31 downto 0);
      conv1402_3925 <= tmp_var; -- 
    end process;
    type_cast_3934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3934_inst_req_0;
      type_cast_3934_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3934_inst_req_1;
      type_cast_3934_inst_ack_1<= rack(0);
      type_cast_3934_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3934_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1272x_x0x_xph_4322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3934_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3938_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3938_inst_req_0;
      type_cast_3938_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3938_inst_req_1;
      type_cast_3938_inst_ack_1<= rack(0);
      type_cast_3938_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3938_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1276x_x1x_xph_4329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3938_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3940_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3940_inst_req_0;
      type_cast_3940_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3940_inst_req_1;
      type_cast_3940_inst_ack_1<= rack(0);
      type_cast_3940_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3940_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul1280_3847,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3940_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3947_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3947_inst_req_0;
      type_cast_3947_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3947_inst_req_1;
      type_cast_3947_inst_ack_1<= rack(0);
      type_cast_3947_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3947_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1327x_x0x_xph_4335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3947_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3952_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3952_inst_req_0;
      type_cast_3952_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3952_inst_req_1;
      type_cast_3952_inst_ack_1<= rack(0);
      type_cast_3952_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3952_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3951_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1333_3953,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3956_inst
    process(conv1333_3953) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1333_3953(31 downto 0);
      type_cast_3956_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3958_inst
    process(conv1335_3880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1335_3880(31 downto 0);
      type_cast_3958_wire <= tmp_var; -- 
    end process;
    type_cast_3973_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3973_inst_req_0;
      type_cast_3973_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3973_inst_req_1;
      type_cast_3973_inst_ack_1<= rack(0);
      type_cast_3973_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3973_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1341_3970,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1342_3974,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3982_inst
    process(conv1333_3953) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1333_3953(31 downto 0);
      type_cast_3982_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3984_inst
    process(add1345_3979) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1345_3979(31 downto 0);
      type_cast_3984_wire <= tmp_var; -- 
    end process;
    type_cast_3997_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3997_inst_req_0;
      type_cast_3997_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3997_inst_req_1;
      type_cast_3997_inst_ack_1<= rack(0);
      type_cast_3997_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3997_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3996_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1350_3998,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4001_inst
    process(conv1350_3998) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1350_3998(31 downto 0);
      type_cast_4001_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4003_inst
    process(conv1335_3880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1335_3880(31 downto 0);
      type_cast_4003_wire <= tmp_var; -- 
    end process;
    type_cast_4018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4018_inst_req_0;
      type_cast_4018_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4018_inst_req_1;
      type_cast_4018_inst_ack_1<= rack(0);
      type_cast_4018_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1358_4015,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1359_4019,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4033_inst
    process(conv1350_3998) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1350_3998(31 downto 0);
      type_cast_4033_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4035_inst
    process(add1363_4030) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1363_4030(31 downto 0);
      type_cast_4035_wire <= tmp_var; -- 
    end process;
    type_cast_4048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4048_inst_req_0;
      type_cast_4048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4048_inst_req_1;
      type_cast_4048_inst_ack_1<= rack(0);
      type_cast_4048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4047_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1370_4049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4053_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4053_inst_req_0;
      type_cast_4053_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4053_inst_req_1;
      type_cast_4053_inst_ack_1<= rack(0);
      type_cast_4053_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4053_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4052_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1374_4054,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4077_inst
    process(add1382_4074) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1382_4074(31 downto 0);
      type_cast_4077_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4082_inst
    process(ASHR_i32_i32_4081_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4081_wire(31 downto 0);
      shr1384_4083 <= tmp_var; -- 
    end process;
    type_cast_4087_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4087_inst_req_0;
      type_cast_4087_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4087_inst_req_1;
      type_cast_4087_inst_ack_1<= rack(0);
      type_cast_4087_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4087_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4086_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1385_4088,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4106_inst_req_0;
      type_cast_4106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4106_inst_req_1;
      type_cast_4106_inst_ack_1<= rack(0);
      type_cast_4106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4105_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1391_4107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4160_inst
    process(add1409_4137) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1409_4137(31 downto 0);
      type_cast_4160_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4165_inst
    process(ASHR_i32_i32_4164_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4164_wire(31 downto 0);
      shr1427_4166 <= tmp_var; -- 
    end process;
    type_cast_4170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4170_inst_req_0;
      type_cast_4170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4170_inst_req_1;
      type_cast_4170_inst_ack_1<= rack(0);
      type_cast_4170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4169_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1428_4171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4185_inst
    process(add1425_4157) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1425_4157(31 downto 0);
      type_cast_4185_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4190_inst
    process(ASHR_i32_i32_4189_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4189_wire(31 downto 0);
      shr1432_4191 <= tmp_var; -- 
    end process;
    type_cast_4195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4195_inst_req_0;
      type_cast_4195_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4195_inst_req_1;
      type_cast_4195_inst_ack_1<= rack(0);
      type_cast_4195_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4195_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4194_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1433_4196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4213_inst_req_0;
      type_cast_4213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4213_inst_req_1;
      type_cast_4213_inst_ack_1<= rack(0);
      type_cast_4213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4212_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1439_4214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4223_inst
    process(add1440_4220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1440_4220(31 downto 0);
      type_cast_4223_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4225_inst
    process(conv1313_3863) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1313_3863(31 downto 0);
      type_cast_4225_wire <= tmp_var; -- 
    end process;
    type_cast_4252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4252_inst_req_0;
      type_cast_4252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4252_inst_req_1;
      type_cast_4252_inst_ack_1<= rack(0);
      type_cast_4252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4251_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1454_4253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4259_inst_req_0;
      type_cast_4259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4259_inst_req_1;
      type_cast_4259_inst_ack_1<= rack(0);
      type_cast_4259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1455_4256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1456_4260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4279_inst_req_0;
      type_cast_4279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4279_inst_req_1;
      type_cast_4279_inst_ack_1<= rack(0);
      type_cast_4279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1462_4276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1467_4280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4296_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4296_inst_req_0;
      type_cast_4296_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4296_inst_req_1;
      type_cast_4296_inst_ack_1<= rack(0);
      type_cast_4296_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4296_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4295_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1470_4297,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4303_inst_req_0;
      type_cast_4303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4303_inst_req_1;
      type_cast_4303_inst_ack_1<= rack(0);
      type_cast_4303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1471_4300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1472_4304,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4325_inst_req_0;
      type_cast_4325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4325_inst_req_1;
      type_cast_4325_inst_ack_1<= rack(0);
      type_cast_4325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1448_4240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4325_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4332_inst_req_0;
      type_cast_4332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4332_inst_req_1;
      type_cast_4332_inst_ack_1<= rack(0);
      type_cast_4332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1276x_x2_3935,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4332_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4334_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4334_inst_req_0;
      type_cast_4334_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4334_inst_req_1;
      type_cast_4334_inst_ack_1<= rack(0);
      type_cast_4334_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4334_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1467x_xi1276x_x2_4285,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4334_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4338_inst_req_0;
      type_cast_4338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4338_inst_req_1;
      type_cast_4338_inst_ack_1<= rack(0);
      type_cast_4338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1327x_x1_3941,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4338_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4340_inst_req_0;
      type_cast_4340_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4340_inst_req_1;
      type_cast_4340_inst_ack_1<= rack(0);
      type_cast_4340_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4340_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1327x_x2_4292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4340_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4347_inst_req_0;
      type_cast_4347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4347_inst_req_1;
      type_cast_4347_inst_ack_1<= rack(0);
      type_cast_4347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1471_4300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4347_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4351_inst_req_0;
      type_cast_4351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4351_inst_req_1;
      type_cast_4351_inst_ack_1<= rack(0);
      type_cast_4351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv1456_4260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4351_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4355_inst_req_0;
      type_cast_4355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4355_inst_req_1;
      type_cast_4355_inst_ack_1<= rack(0);
      type_cast_4355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1455_4256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4355_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4359_inst_req_0;
      type_cast_4359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4359_inst_req_1;
      type_cast_4359_inst_ack_1<= rack(0);
      type_cast_4359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1455x_xlcssa_4352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1493_4360,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4369_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4369_inst_req_0;
      type_cast_4369_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4369_inst_req_1;
      type_cast_4369_inst_ack_1<= rack(0);
      type_cast_4369_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4369_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1471x_xlcssa_4344,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1499_4370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4397_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4397_inst_req_0;
      type_cast_4397_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4397_inst_req_1;
      type_cast_4397_inst_ack_1<= rack(0);
      type_cast_4397_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4397_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1509_4388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1534_4398,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4401_inst_req_0;
      type_cast_4401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4401_inst_req_1;
      type_cast_4401_inst_ack_1<= rack(0);
      type_cast_4401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1521_4391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1542_4402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4405_inst_req_0;
      type_cast_4405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4405_inst_req_1;
      type_cast_4405_inst_ack_1<= rack(0);
      type_cast_4405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1525_4394,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1544_4406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4414_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4414_inst_req_0;
      type_cast_4414_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4414_inst_req_1;
      type_cast_4414_inst_ack_1<= rack(0);
      type_cast_4414_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4414_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1505_4385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1556_4415,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4418_inst_req_0;
      type_cast_4418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4418_inst_req_1;
      type_cast_4418_inst_ack_1<= rack(0);
      type_cast_4418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1521_4391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1592_4419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4428_inst
    process(sext1753_4425) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1753_4425(31 downto 0);
      type_cast_4428_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4433_inst
    process(ASHR_i32_i32_4432_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4432_wire(31 downto 0);
      conv1598_4434 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4454_inst
    process(sext1713_4451) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1713_4451(31 downto 0);
      type_cast_4454_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4459_inst
    process(ASHR_i32_i32_4458_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4458_wire(31 downto 0);
      conv1622_4460 <= tmp_var; -- 
    end process;
    type_cast_4469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4469_inst_req_0;
      type_cast_4469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4469_inst_req_1;
      type_cast_4469_inst_ack_1<= rack(0);
      type_cast_4469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1489x_x0x_xph_4843,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4469_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4473_inst_req_0;
      type_cast_4473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4473_inst_req_1;
      type_cast_4473_inst_ack_1<= rack(0);
      type_cast_4473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1501_4382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4473_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4475_inst_req_0;
      type_cast_4475_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4475_inst_req_1;
      type_cast_4475_inst_ack_1<= rack(0);
      type_cast_4475_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1497x_x1x_xph_4850,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4475_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4479_inst_req_0;
      type_cast_4479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4479_inst_req_1;
      type_cast_4479_inst_ack_1<= rack(0);
      type_cast_4479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1494_4366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4479_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4481_inst_req_0;
      type_cast_4481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4481_inst_req_1;
      type_cast_4481_inst_ack_1<= rack(0);
      type_cast_4481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1548x_x0x_xph_4856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4481_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4486_inst_req_0;
      type_cast_4486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4486_inst_req_1;
      type_cast_4486_inst_ack_1<= rack(0);
      type_cast_4486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4485_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1554_4487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4490_inst
    process(conv1554_4487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1554_4487(31 downto 0);
      type_cast_4490_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4492_inst
    process(conv1556_4415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1556_4415(31 downto 0);
      type_cast_4492_wire <= tmp_var; -- 
    end process;
    type_cast_4507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4507_inst_req_0;
      type_cast_4507_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4507_inst_req_1;
      type_cast_4507_inst_ack_1<= rack(0);
      type_cast_4507_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4507_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1562_4504,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1563_4508,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4516_inst
    process(conv1554_4487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1554_4487(31 downto 0);
      type_cast_4516_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4518_inst
    process(add1566_4513) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1566_4513(31 downto 0);
      type_cast_4518_wire <= tmp_var; -- 
    end process;
    type_cast_4531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4531_inst_req_0;
      type_cast_4531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4531_inst_req_1;
      type_cast_4531_inst_ack_1<= rack(0);
      type_cast_4531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4530_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1571_4532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4535_inst
    process(conv1571_4532) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1571_4532(31 downto 0);
      type_cast_4535_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4537_inst
    process(conv1556_4415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1556_4415(31 downto 0);
      type_cast_4537_wire <= tmp_var; -- 
    end process;
    type_cast_4552_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4552_inst_req_0;
      type_cast_4552_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4552_inst_req_1;
      type_cast_4552_inst_ack_1<= rack(0);
      type_cast_4552_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4552_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1579_4549,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1580_4553,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4561_inst
    process(conv1571_4532) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1571_4532(31 downto 0);
      type_cast_4561_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4563_inst
    process(add1583_4558) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1583_4558(31 downto 0);
      type_cast_4563_wire <= tmp_var; -- 
    end process;
    type_cast_4576_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4576_inst_req_0;
      type_cast_4576_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4576_inst_req_1;
      type_cast_4576_inst_ack_1<= rack(0);
      type_cast_4576_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4576_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4575_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1590_4577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4581_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4581_inst_req_0;
      type_cast_4581_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4581_inst_req_1;
      type_cast_4581_inst_ack_1<= rack(0);
      type_cast_4581_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4581_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4580_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1594_4582,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4605_inst
    process(add1602_4602) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1602_4602(31 downto 0);
      type_cast_4605_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4610_inst
    process(ASHR_i32_i32_4609_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4609_wire(31 downto 0);
      shr1604_4611 <= tmp_var; -- 
    end process;
    type_cast_4615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4615_inst_req_0;
      type_cast_4615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4615_inst_req_1;
      type_cast_4615_inst_ack_1<= rack(0);
      type_cast_4615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4614_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1605_4616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4634_inst_req_0;
      type_cast_4634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4634_inst_req_1;
      type_cast_4634_inst_ack_1<= rack(0);
      type_cast_4634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4633_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1611_4635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4688_inst
    process(add1629_4665) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1629_4665(31 downto 0);
      type_cast_4688_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4693_inst
    process(ASHR_i32_i32_4692_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4692_wire(31 downto 0);
      shr1647_4694 <= tmp_var; -- 
    end process;
    type_cast_4698_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4698_inst_req_0;
      type_cast_4698_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4698_inst_req_1;
      type_cast_4698_inst_ack_1<= rack(0);
      type_cast_4698_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4698_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4697_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1648_4699,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4713_inst
    process(add1645_4685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1645_4685(31 downto 0);
      type_cast_4713_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4718_inst
    process(ASHR_i32_i32_4717_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4717_wire(31 downto 0);
      shr1652_4719 <= tmp_var; -- 
    end process;
    type_cast_4723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4723_inst_req_0;
      type_cast_4723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4723_inst_req_1;
      type_cast_4723_inst_ack_1<= rack(0);
      type_cast_4723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4722_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1653_4724,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4741_inst_req_0;
      type_cast_4741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4741_inst_req_1;
      type_cast_4741_inst_ack_1<= rack(0);
      type_cast_4741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4740_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1659_4742,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4751_inst
    process(add1660_4748) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1660_4748(31 downto 0);
      type_cast_4751_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4753_inst
    process(conv1534_4398) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1534_4398(31 downto 0);
      type_cast_4753_wire <= tmp_var; -- 
    end process;
    type_cast_4780_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4780_inst_req_0;
      type_cast_4780_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4780_inst_req_1;
      type_cast_4780_inst_ack_1<= rack(0);
      type_cast_4780_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4780_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4779_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1674_4781,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4787_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4787_inst_req_0;
      type_cast_4787_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4787_inst_req_1;
      type_cast_4787_inst_ack_1<= rack(0);
      type_cast_4787_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4787_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1675_4784,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1676_4788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4801_inst_req_0;
      type_cast_4801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4801_inst_req_1;
      type_cast_4801_inst_ack_1<= rack(0);
      type_cast_4801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1681_4798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1686_4802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4817_inst_req_0;
      type_cast_4817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4817_inst_req_1;
      type_cast_4817_inst_ack_1<= rack(0);
      type_cast_4817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4816_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1689_4818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4824_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4824_inst_req_0;
      type_cast_4824_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4824_inst_req_1;
      type_cast_4824_inst_ack_1<= rack(0);
      type_cast_4824_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4824_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1690_4821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1691_4825,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4849_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4849_inst_req_0;
      type_cast_4849_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4849_inst_req_1;
      type_cast_4849_inst_ack_1<= rack(0);
      type_cast_4849_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4849_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1668_4768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4849_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4853_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4853_inst_req_0;
      type_cast_4853_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4853_inst_req_1;
      type_cast_4853_inst_ack_1<= rack(0);
      type_cast_4853_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4853_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1497x_x2_4470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4853_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4855_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4855_inst_req_0;
      type_cast_4855_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4855_inst_req_1;
      type_cast_4855_inst_ack_1<= rack(0);
      type_cast_4855_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4855_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1686x_xi1497x_x2_4807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4855_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4859_inst_req_0;
      type_cast_4859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4859_inst_req_1;
      type_cast_4859_inst_ack_1<= rack(0);
      type_cast_4859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1548x_x1_4476,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4859_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4861_inst_req_0;
      type_cast_4861_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4861_inst_req_1;
      type_cast_4861_inst_ack_1<= rack(0);
      type_cast_4861_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4861_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1548x_x2_4813,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4861_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_676_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_676_inst_req_0;
      type_cast_676_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_676_inst_req_1;
      type_cast_676_inst_ack_1<= rack(0);
      type_cast_676_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_676_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp2_664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv21_677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_680_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_680_inst_req_0;
      type_cast_680_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_680_inst_req_1;
      type_cast_680_inst_ack_1<= rack(0);
      type_cast_680_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_680_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_667,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_681,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_684_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_684_inst_req_0;
      type_cast_684_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_684_inst_req_1;
      type_cast_684_inst_ack_1<= rack(0);
      type_cast_684_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_684_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_685,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_688_inst_req_0;
      type_cast_688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_688_inst_req_1;
      type_cast_688_inst_ack_1<= rack(0);
      type_cast_688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_697_inst_req_0;
      type_cast_697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_697_inst_req_1;
      type_cast_697_inst_ack_1<= rack(0);
      type_cast_697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_701_inst_req_0;
      type_cast_701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_701_inst_req_1;
      type_cast_701_inst_ack_1<= rack(0);
      type_cast_701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_712_inst
    process(sext1746_708) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1746_708(31 downto 0);
      type_cast_712_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_717_inst
    process(ASHR_i32_i32_716_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_716_wire(31 downto 0);
      conv76_718 <= tmp_var; -- 
    end process;
    -- interlock type_cast_738_inst
    process(sext_735) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_735(31 downto 0);
      type_cast_738_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_743_inst
    process(ASHR_i32_i32_742_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_742_wire(31 downto 0);
      conv94_744 <= tmp_var; -- 
    end process;
    type_cast_753_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_753_inst_req_0;
      type_cast_753_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_753_inst_req_1;
      type_cast_753_inst_ack_1<= rack(0);
      type_cast_753_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_753_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_1155,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_753_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_760_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_760_inst_req_0;
      type_cast_760_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_760_inst_req_1;
      type_cast_760_inst_ack_1<= rack(0);
      type_cast_760_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_760_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_1161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_760_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_767_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_767_inst_req_0;
      type_cast_767_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_767_inst_req_1;
      type_cast_767_inst_ack_1<= rack(0);
      type_cast_767_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_767_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_1167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_767_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_772_inst_req_0;
      type_cast_772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_772_inst_req_1;
      type_cast_772_inst_ack_1<= rack(0);
      type_cast_772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_771_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_776_inst
    process(conv36_773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv36_773(31 downto 0);
      type_cast_776_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_778_inst
    process(conv38_698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv38_698(31 downto 0);
      type_cast_778_wire <= tmp_var; -- 
    end process;
    type_cast_793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_793_inst_req_0;
      type_cast_793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_793_inst_req_1;
      type_cast_793_inst_ack_1<= rack(0);
      type_cast_793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp42_790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_808_inst
    process(conv36_773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv36_773(31 downto 0);
      type_cast_808_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_810_inst
    process(add_805) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_805(31 downto 0);
      type_cast_810_wire <= tmp_var; -- 
    end process;
    type_cast_823_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_823_inst_req_0;
      type_cast_823_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_823_inst_req_1;
      type_cast_823_inst_ack_1<= rack(0);
      type_cast_823_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_823_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_822_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_824,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_827_inst
    process(conv50_824) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv50_824(31 downto 0);
      type_cast_827_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_829_inst
    process(conv38_698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv38_698(31 downto 0);
      type_cast_829_wire <= tmp_var; -- 
    end process;
    type_cast_844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_844_inst_req_0;
      type_cast_844_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_844_inst_req_1;
      type_cast_844_inst_ack_1<= rack(0);
      type_cast_844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp58_841,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_845,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_859_inst
    process(conv50_824) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv50_824(31 downto 0);
      type_cast_859_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_861_inst
    process(add63_856) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add63_856(31 downto 0);
      type_cast_861_wire <= tmp_var; -- 
    end process;
    type_cast_874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_874_inst_req_0;
      type_cast_874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_874_inst_req_1;
      type_cast_874_inst_ack_1<= rack(0);
      type_cast_874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_873_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_879_inst_req_0;
      type_cast_879_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_879_inst_req_1;
      type_cast_879_inst_ack_1<= rack(0);
      type_cast_879_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_879_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_878_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_880,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_903_inst
    process(add80_900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add80_900(31 downto 0);
      type_cast_903_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_908_inst
    process(ASHR_i32_i32_907_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_907_wire(31 downto 0);
      shr_909 <= tmp_var; -- 
    end process;
    type_cast_914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_914_inst_req_0;
      type_cast_914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_914_inst_req_1;
      type_cast_914_inst_ack_1<= rack(0);
      type_cast_914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_913_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_933_inst_req_0;
      type_cast_933_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_933_inst_req_1;
      type_cast_933_inst_ack_1<= rack(0);
      type_cast_933_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_932_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_987_inst
    process(add101_964) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add101_964(31 downto 0);
      type_cast_987_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_992_inst
    process(ASHR_i32_i32_991_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_991_wire(31 downto 0);
      shr119_993 <= tmp_var; -- 
    end process;
    type_cast_997_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_997_inst_req_0;
      type_cast_997_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_997_inst_req_1;
      type_cast_997_inst_ack_1<= rack(0);
      type_cast_997_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_997_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_996_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom120_998,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_col_high_1082_gather_scatter
    process(LOAD_col_high_1082_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1082_data_0;
      ov(7 downto 0) := iv;
      tmp144_1083 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1368_gather_scatter
    process(LOAD_col_high_1368_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1368_data_0;
      ov(7 downto 0) := iv;
      tmp262_1369 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1603_gather_scatter
    process(LOAD_col_high_1603_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1603_data_0;
      ov(7 downto 0) := iv;
      tmp358_1604 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1882_gather_scatter
    process(LOAD_col_high_1882_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1882_data_0;
      ov(7 downto 0) := iv;
      tmp478_1883 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2123_gather_scatter
    process(LOAD_col_high_2123_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2123_data_0;
      ov(7 downto 0) := iv;
      tmp575_2124 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2422_gather_scatter
    process(LOAD_col_high_2422_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2422_data_0;
      ov(7 downto 0) := iv;
      tmp700_2423 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2657_gather_scatter
    process(LOAD_col_high_2657_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2657_data_0;
      ov(7 downto 0) := iv;
      tmp796_2658 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2942_gather_scatter
    process(LOAD_col_high_2942_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2942_data_0;
      ov(7 downto 0) := iv;
      tmp917_2943 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3183_gather_scatter
    process(LOAD_col_high_3183_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3183_data_0;
      ov(7 downto 0) := iv;
      tmp1014_3184 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3494_gather_scatter
    process(LOAD_col_high_3494_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3494_data_0;
      ov(7 downto 0) := iv;
      tmp1141_3495 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3729_gather_scatter
    process(LOAD_col_high_3729_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3729_data_0;
      ov(7 downto 0) := iv;
      tmp1237_3730 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4014_gather_scatter
    process(LOAD_col_high_4014_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4014_data_0;
      ov(7 downto 0) := iv;
      tmp1358_4015 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4255_gather_scatter
    process(LOAD_col_high_4255_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4255_data_0;
      ov(7 downto 0) := iv;
      tmp1455_4256 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4548_gather_scatter
    process(LOAD_col_high_4548_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4548_data_0;
      ov(7 downto 0) := iv;
      tmp1579_4549 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4783_gather_scatter
    process(LOAD_col_high_4783_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4783_data_0;
      ov(7 downto 0) := iv;
      tmp1675_4784 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_666_gather_scatter
    process(LOAD_col_high_666_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_666_data_0;
      ov(7 downto 0) := iv;
      tmp5_667 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_840_gather_scatter
    process(LOAD_col_high_840_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_840_data_0;
      ov(7 downto 0) := iv;
      tmp58_841 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_1200_gather_scatter
    process(LOAD_depth_high_1200_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_1200_data_0;
      ov(7 downto 0) := iv;
      tmp191_1201 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_1714_gather_scatter
    process(LOAD_depth_high_1714_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_1714_data_0;
      ov(7 downto 0) := iv;
      tmp407_1715 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_2255_gather_scatter
    process(LOAD_depth_high_2255_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_2255_data_0;
      ov(7 downto 0) := iv;
      tmp629_2256 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_2768_gather_scatter
    process(LOAD_depth_high_2768_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_2768_data_0;
      ov(7 downto 0) := iv;
      tmp845_2769 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_3321_gather_scatter
    process(LOAD_depth_high_3321_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_3321_data_0;
      ov(7 downto 0) := iv;
      tmp1069_3322 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_3852_gather_scatter
    process(LOAD_depth_high_3852_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_3852_data_0;
      ov(7 downto 0) := iv;
      tmp1288_3853 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_4387_gather_scatter
    process(LOAD_depth_high_4387_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_4387_data_0;
      ov(7 downto 0) := iv;
      tmp1509_4388 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_663_gather_scatter
    process(LOAD_depth_high_663_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_663_data_0;
      ov(7 downto 0) := iv;
      tmp2_664 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_col_high_1206_gather_scatter
    process(LOAD_out_col_high_1206_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_1206_data_0;
      ov(7 downto 0) := iv;
      tmp207_1207 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_col_high_1720_gather_scatter
    process(LOAD_out_col_high_1720_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_1720_data_0;
      ov(7 downto 0) := iv;
      tmp423_1721 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_col_high_2261_gather_scatter
    process(LOAD_out_col_high_2261_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_2261_data_0;
      ov(7 downto 0) := iv;
      tmp645_2262 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_col_high_2774_gather_scatter
    process(LOAD_out_col_high_2774_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_2774_data_0;
      ov(7 downto 0) := iv;
      tmp861_2775 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_col_high_3327_gather_scatter
    process(LOAD_out_col_high_3327_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_3327_data_0;
      ov(7 downto 0) := iv;
      tmp1085_3328 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_col_high_3858_gather_scatter
    process(LOAD_out_col_high_3858_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_3858_data_0;
      ov(7 downto 0) := iv;
      tmp1304_3859 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_col_high_4393_gather_scatter
    process(LOAD_out_col_high_4393_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_4393_data_0;
      ov(7 downto 0) := iv;
      tmp1525_4394 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_col_high_672_gather_scatter
    process(LOAD_out_col_high_672_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_col_high_672_data_0;
      ov(7 downto 0) := iv;
      tmp14_673 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_1203_gather_scatter
    process(LOAD_out_depth_high_1203_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_1203_data_0;
      ov(7 downto 0) := iv;
      tmp203_1204 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_1717_gather_scatter
    process(LOAD_out_depth_high_1717_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_1717_data_0;
      ov(7 downto 0) := iv;
      tmp419_1718 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_2258_gather_scatter
    process(LOAD_out_depth_high_2258_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_2258_data_0;
      ov(7 downto 0) := iv;
      tmp641_2259 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_2771_gather_scatter
    process(LOAD_out_depth_high_2771_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_2771_data_0;
      ov(7 downto 0) := iv;
      tmp857_2772 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_3324_gather_scatter
    process(LOAD_out_depth_high_3324_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_3324_data_0;
      ov(7 downto 0) := iv;
      tmp1081_3325 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_3855_gather_scatter
    process(LOAD_out_depth_high_3855_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_3855_data_0;
      ov(7 downto 0) := iv;
      tmp1300_3856 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_4390_gather_scatter
    process(LOAD_out_depth_high_4390_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_4390_data_0;
      ov(7 downto 0) := iv;
      tmp1521_4391 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_out_depth_high_669_gather_scatter
    process(LOAD_out_depth_high_669_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_out_depth_high_669_data_0;
      ov(7 downto 0) := iv;
      tmp11_670 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_1197_gather_scatter
    process(LOAD_pad_1197_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1197_data_0;
      ov(7 downto 0) := iv;
      tmp187_1198 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_1711_gather_scatter
    process(LOAD_pad_1711_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1711_data_0;
      ov(7 downto 0) := iv;
      tmp403_1712 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_2252_gather_scatter
    process(LOAD_pad_2252_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_2252_data_0;
      ov(7 downto 0) := iv;
      tmp625_2253 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_2765_gather_scatter
    process(LOAD_pad_2765_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_2765_data_0;
      ov(7 downto 0) := iv;
      tmp841_2766 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_3318_gather_scatter
    process(LOAD_pad_3318_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_3318_data_0;
      ov(7 downto 0) := iv;
      tmp1065_3319 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_3849_gather_scatter
    process(LOAD_pad_3849_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_3849_data_0;
      ov(7 downto 0) := iv;
      tmp1284_3850 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_4384_gather_scatter
    process(LOAD_pad_4384_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_4384_data_0;
      ov(7 downto 0) := iv;
      tmp1505_4385 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_660_gather_scatter
    process(LOAD_pad_660_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_660_data_0;
      ov(7 downto 0) := iv;
      tmp_661 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1126_gather_scatter
    process(LOAD_row_high_1126_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1126_data_0;
      ov(7 downto 0) := iv;
      tmp159_1127 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1317_gather_scatter
    process(LOAD_row_high_1317_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1317_data_0;
      ov(7 downto 0) := iv;
      tmp244_1318 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1640_gather_scatter
    process(LOAD_row_high_1640_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1640_data_0;
      ov(7 downto 0) := iv;
      tmp373_1641 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1831_gather_scatter
    process(LOAD_row_high_1831_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1831_data_0;
      ov(7 downto 0) := iv;
      tmp460_1832 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2167_gather_scatter
    process(LOAD_row_high_2167_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2167_data_0;
      ov(7 downto 0) := iv;
      tmp591_2168 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2371_gather_scatter
    process(LOAD_row_high_2371_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2371_data_0;
      ov(7 downto 0) := iv;
      tmp682_2372 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2694_gather_scatter
    process(LOAD_row_high_2694_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2694_data_0;
      ov(7 downto 0) := iv;
      tmp811_2695 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2885_gather_scatter
    process(LOAD_row_high_2885_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2885_data_0;
      ov(7 downto 0) := iv;
      tmp898_2886 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3227_gather_scatter
    process(LOAD_row_high_3227_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3227_data_0;
      ov(7 downto 0) := iv;
      tmp1030_3228 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3437_gather_scatter
    process(LOAD_row_high_3437_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3437_data_0;
      ov(7 downto 0) := iv;
      tmp1122_3438 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3766_gather_scatter
    process(LOAD_row_high_3766_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3766_data_0;
      ov(7 downto 0) := iv;
      tmp1252_3767 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3969_gather_scatter
    process(LOAD_row_high_3969_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3969_data_0;
      ov(7 downto 0) := iv;
      tmp1341_3970 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4299_gather_scatter
    process(LOAD_row_high_4299_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4299_data_0;
      ov(7 downto 0) := iv;
      tmp1471_4300 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4503_gather_scatter
    process(LOAD_row_high_4503_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4503_data_0;
      ov(7 downto 0) := iv;
      tmp1562_4504 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4820_gather_scatter
    process(LOAD_row_high_4820_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4820_data_0;
      ov(7 downto 0) := iv;
      tmp1690_4821 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_789_gather_scatter
    process(LOAD_row_high_789_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_789_data_0;
      ov(7 downto 0) := iv;
      tmp42_790 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1003_index_1_rename
    process(R_idxprom120_1002_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom120_1002_resized;
      ov(13 downto 0) := iv;
      R_idxprom120_1002_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1003_index_1_resize
    process(idxprom120_998) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom120_998;
      ov := iv(13 downto 0);
      R_idxprom120_1002_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1003_root_address_inst
    process(array_obj_ref_1003_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1003_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1003_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1028_index_1_rename
    process(R_idxprom125_1027_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom125_1027_resized;
      ov(13 downto 0) := iv;
      R_idxprom125_1027_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1028_index_1_resize
    process(idxprom125_1023) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom125_1023;
      ov := iv(13 downto 0);
      R_idxprom125_1027_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1028_root_address_inst
    process(array_obj_ref_1028_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1028_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1028_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_index_1_rename
    process(R_idxprom288_1440_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom288_1440_resized;
      ov(13 downto 0) := iv;
      R_idxprom288_1440_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_index_1_resize
    process(idxprom288_1436) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom288_1436;
      ov := iv(13 downto 0);
      R_idxprom288_1440_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1441_root_address_inst
    process(array_obj_ref_1441_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1441_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1441_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1524_index_1_rename
    process(R_idxprom331_1523_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom331_1523_resized;
      ov(13 downto 0) := iv;
      R_idxprom331_1523_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1524_index_1_resize
    process(idxprom331_1519) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom331_1519;
      ov := iv(13 downto 0);
      R_idxprom331_1523_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1524_root_address_inst
    process(array_obj_ref_1524_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1524_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1524_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1549_index_1_rename
    process(R_idxprom336_1548_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom336_1548_resized;
      ov(13 downto 0) := iv;
      R_idxprom336_1548_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1549_index_1_resize
    process(idxprom336_1544) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom336_1544;
      ov := iv(13 downto 0);
      R_idxprom336_1548_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1549_root_address_inst
    process(array_obj_ref_1549_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1549_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1549_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1961_index_1_rename
    process(R_idxprom505_1960_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom505_1960_resized;
      ov(13 downto 0) := iv;
      R_idxprom505_1960_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1961_index_1_resize
    process(idxprom505_1956) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom505_1956;
      ov := iv(13 downto 0);
      R_idxprom505_1960_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1961_root_address_inst
    process(array_obj_ref_1961_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1961_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1961_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2044_index_1_rename
    process(R_idxprom548_2043_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom548_2043_resized;
      ov(13 downto 0) := iv;
      R_idxprom548_2043_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2044_index_1_resize
    process(idxprom548_2039) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom548_2039;
      ov := iv(13 downto 0);
      R_idxprom548_2043_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2044_root_address_inst
    process(array_obj_ref_2044_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2044_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2044_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2069_index_1_rename
    process(R_idxprom553_2068_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom553_2068_resized;
      ov(13 downto 0) := iv;
      R_idxprom553_2068_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2069_index_1_resize
    process(idxprom553_2064) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom553_2064;
      ov := iv(13 downto 0);
      R_idxprom553_2068_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2069_root_address_inst
    process(array_obj_ref_2069_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2069_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2069_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2495_index_1_rename
    process(R_idxprom726_2494_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom726_2494_resized;
      ov(13 downto 0) := iv;
      R_idxprom726_2494_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2495_index_1_resize
    process(idxprom726_2490) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom726_2490;
      ov := iv(13 downto 0);
      R_idxprom726_2494_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2495_root_address_inst
    process(array_obj_ref_2495_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2495_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2495_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2578_index_1_rename
    process(R_idxprom769_2577_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom769_2577_resized;
      ov(13 downto 0) := iv;
      R_idxprom769_2577_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2578_index_1_resize
    process(idxprom769_2573) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom769_2573;
      ov := iv(13 downto 0);
      R_idxprom769_2577_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2578_root_address_inst
    process(array_obj_ref_2578_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2578_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2578_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2603_index_1_rename
    process(R_idxprom774_2602_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom774_2602_resized;
      ov(13 downto 0) := iv;
      R_idxprom774_2602_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2603_index_1_resize
    process(idxprom774_2598) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom774_2598;
      ov := iv(13 downto 0);
      R_idxprom774_2602_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2603_root_address_inst
    process(array_obj_ref_2603_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2603_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2603_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3021_index_1_rename
    process(R_idxprom944_3020_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom944_3020_resized;
      ov(13 downto 0) := iv;
      R_idxprom944_3020_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3021_index_1_resize
    process(idxprom944_3016) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom944_3016;
      ov := iv(13 downto 0);
      R_idxprom944_3020_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3021_root_address_inst
    process(array_obj_ref_3021_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3021_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3021_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3104_index_1_rename
    process(R_idxprom987_3103_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom987_3103_resized;
      ov(13 downto 0) := iv;
      R_idxprom987_3103_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3104_index_1_resize
    process(idxprom987_3099) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom987_3099;
      ov := iv(13 downto 0);
      R_idxprom987_3103_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3104_root_address_inst
    process(array_obj_ref_3104_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3104_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3104_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3129_index_1_rename
    process(R_idxprom992_3128_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom992_3128_resized;
      ov(13 downto 0) := iv;
      R_idxprom992_3128_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3129_index_1_resize
    process(idxprom992_3124) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom992_3124;
      ov := iv(13 downto 0);
      R_idxprom992_3128_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3129_root_address_inst
    process(array_obj_ref_3129_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3129_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3129_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3567_index_1_rename
    process(R_idxprom1167_3566_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1167_3566_resized;
      ov(13 downto 0) := iv;
      R_idxprom1167_3566_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3567_index_1_resize
    process(idxprom1167_3562) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1167_3562;
      ov := iv(13 downto 0);
      R_idxprom1167_3566_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3567_root_address_inst
    process(array_obj_ref_3567_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3567_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3567_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3650_index_1_rename
    process(R_idxprom1210_3649_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1210_3649_resized;
      ov(13 downto 0) := iv;
      R_idxprom1210_3649_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3650_index_1_resize
    process(idxprom1210_3645) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1210_3645;
      ov := iv(13 downto 0);
      R_idxprom1210_3649_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3650_root_address_inst
    process(array_obj_ref_3650_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3650_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3650_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3675_index_1_rename
    process(R_idxprom1215_3674_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1215_3674_resized;
      ov(13 downto 0) := iv;
      R_idxprom1215_3674_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3675_index_1_resize
    process(idxprom1215_3670) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1215_3670;
      ov := iv(13 downto 0);
      R_idxprom1215_3674_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3675_root_address_inst
    process(array_obj_ref_3675_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3675_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3675_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4093_index_1_rename
    process(R_idxprom1385_4092_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1385_4092_resized;
      ov(13 downto 0) := iv;
      R_idxprom1385_4092_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4093_index_1_resize
    process(idxprom1385_4088) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1385_4088;
      ov := iv(13 downto 0);
      R_idxprom1385_4092_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4093_root_address_inst
    process(array_obj_ref_4093_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4093_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4093_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4176_index_1_rename
    process(R_idxprom1428_4175_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1428_4175_resized;
      ov(13 downto 0) := iv;
      R_idxprom1428_4175_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4176_index_1_resize
    process(idxprom1428_4171) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1428_4171;
      ov := iv(13 downto 0);
      R_idxprom1428_4175_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4176_root_address_inst
    process(array_obj_ref_4176_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4176_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4176_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4201_index_1_rename
    process(R_idxprom1433_4200_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1433_4200_resized;
      ov(13 downto 0) := iv;
      R_idxprom1433_4200_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4201_index_1_resize
    process(idxprom1433_4196) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1433_4196;
      ov := iv(13 downto 0);
      R_idxprom1433_4200_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4201_root_address_inst
    process(array_obj_ref_4201_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4201_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4201_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4621_index_1_rename
    process(R_idxprom1605_4620_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1605_4620_resized;
      ov(13 downto 0) := iv;
      R_idxprom1605_4620_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4621_index_1_resize
    process(idxprom1605_4616) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1605_4616;
      ov := iv(13 downto 0);
      R_idxprom1605_4620_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4621_root_address_inst
    process(array_obj_ref_4621_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4621_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4621_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4704_index_1_rename
    process(R_idxprom1648_4703_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1648_4703_resized;
      ov(13 downto 0) := iv;
      R_idxprom1648_4703_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4704_index_1_resize
    process(idxprom1648_4699) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1648_4699;
      ov := iv(13 downto 0);
      R_idxprom1648_4703_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4704_root_address_inst
    process(array_obj_ref_4704_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4704_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4704_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4729_index_1_rename
    process(R_idxprom1653_4728_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1653_4728_resized;
      ov(13 downto 0) := iv;
      R_idxprom1653_4728_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4729_index_1_resize
    process(idxprom1653_4724) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1653_4724;
      ov := iv(13 downto 0);
      R_idxprom1653_4728_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4729_root_address_inst
    process(array_obj_ref_4729_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4729_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4729_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_920_index_1_rename
    process(R_idxprom_919_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_919_resized;
      ov(13 downto 0) := iv;
      R_idxprom_919_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_920_index_1_resize
    process(idxprom_915) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_915;
      ov := iv(13 downto 0);
      R_idxprom_919_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_920_root_address_inst
    process(array_obj_ref_920_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_920_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_920_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1008_addr_0
    process(ptr_deref_1008_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1008_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1008_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1008_base_resize
    process(arrayidx121_1005) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx121_1005;
      ov := iv(13 downto 0);
      ptr_deref_1008_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1008_gather_scatter
    process(ptr_deref_1008_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1008_data_0;
      ov(63 downto 0) := iv;
      tmp122_1009 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1008_root_address_inst
    process(ptr_deref_1008_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1008_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1008_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1032_addr_0
    process(ptr_deref_1032_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1032_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1032_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1032_base_resize
    process(arrayidx126_1030) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx126_1030;
      ov := iv(13 downto 0);
      ptr_deref_1032_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1032_gather_scatter
    process(tmp122_1009) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp122_1009;
      ov(63 downto 0) := iv;
      ptr_deref_1032_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1032_root_address_inst
    process(ptr_deref_1032_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1032_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1032_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1445_addr_0
    process(ptr_deref_1445_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1445_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1445_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1445_base_resize
    process(arrayidx289_1443) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx289_1443;
      ov := iv(13 downto 0);
      ptr_deref_1445_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1445_gather_scatter
    process(type_cast_1447_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1447_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1445_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1445_root_address_inst
    process(ptr_deref_1445_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1445_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1445_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1529_addr_0
    process(ptr_deref_1529_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1529_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1529_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1529_base_resize
    process(arrayidx332_1526) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx332_1526;
      ov := iv(13 downto 0);
      ptr_deref_1529_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1529_gather_scatter
    process(ptr_deref_1529_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1529_data_0;
      ov(63 downto 0) := iv;
      tmp333_1530 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1529_root_address_inst
    process(ptr_deref_1529_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1529_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1529_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1553_addr_0
    process(ptr_deref_1553_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1553_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1553_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1553_base_resize
    process(arrayidx337_1551) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx337_1551;
      ov := iv(13 downto 0);
      ptr_deref_1553_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1553_gather_scatter
    process(tmp333_1530) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp333_1530;
      ov(63 downto 0) := iv;
      ptr_deref_1553_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1553_root_address_inst
    process(ptr_deref_1553_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1553_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1553_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1965_addr_0
    process(ptr_deref_1965_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1965_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1965_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1965_base_resize
    process(arrayidx506_1963) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx506_1963;
      ov := iv(13 downto 0);
      ptr_deref_1965_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1965_gather_scatter
    process(type_cast_1967_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1967_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1965_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1965_root_address_inst
    process(ptr_deref_1965_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1965_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1965_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2049_addr_0
    process(ptr_deref_2049_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2049_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2049_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2049_base_resize
    process(arrayidx549_2046) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx549_2046;
      ov := iv(13 downto 0);
      ptr_deref_2049_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2049_gather_scatter
    process(ptr_deref_2049_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2049_data_0;
      ov(63 downto 0) := iv;
      tmp550_2050 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2049_root_address_inst
    process(ptr_deref_2049_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2049_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2049_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_addr_0
    process(ptr_deref_2073_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2073_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2073_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_base_resize
    process(arrayidx554_2071) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx554_2071;
      ov := iv(13 downto 0);
      ptr_deref_2073_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_gather_scatter
    process(tmp550_2050) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp550_2050;
      ov(63 downto 0) := iv;
      ptr_deref_2073_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_root_address_inst
    process(ptr_deref_2073_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2073_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2073_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2499_addr_0
    process(ptr_deref_2499_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2499_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2499_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2499_base_resize
    process(arrayidx727_2497) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx727_2497;
      ov := iv(13 downto 0);
      ptr_deref_2499_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2499_gather_scatter
    process(type_cast_2501_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2501_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2499_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2499_root_address_inst
    process(ptr_deref_2499_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2499_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2499_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2583_addr_0
    process(ptr_deref_2583_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2583_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2583_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2583_base_resize
    process(arrayidx770_2580) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx770_2580;
      ov := iv(13 downto 0);
      ptr_deref_2583_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2583_gather_scatter
    process(ptr_deref_2583_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2583_data_0;
      ov(63 downto 0) := iv;
      tmp771_2584 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2583_root_address_inst
    process(ptr_deref_2583_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2583_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2583_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2607_addr_0
    process(ptr_deref_2607_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2607_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2607_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2607_base_resize
    process(arrayidx775_2605) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx775_2605;
      ov := iv(13 downto 0);
      ptr_deref_2607_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2607_gather_scatter
    process(tmp771_2584) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp771_2584;
      ov(63 downto 0) := iv;
      ptr_deref_2607_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2607_root_address_inst
    process(ptr_deref_2607_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2607_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2607_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3025_addr_0
    process(ptr_deref_3025_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3025_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3025_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3025_base_resize
    process(arrayidx945_3023) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx945_3023;
      ov := iv(13 downto 0);
      ptr_deref_3025_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3025_gather_scatter
    process(type_cast_3027_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3027_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3025_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3025_root_address_inst
    process(ptr_deref_3025_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3025_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3025_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3109_addr_0
    process(ptr_deref_3109_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3109_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3109_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3109_base_resize
    process(arrayidx988_3106) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx988_3106;
      ov := iv(13 downto 0);
      ptr_deref_3109_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3109_gather_scatter
    process(ptr_deref_3109_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3109_data_0;
      ov(63 downto 0) := iv;
      tmp989_3110 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3109_root_address_inst
    process(ptr_deref_3109_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3109_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3109_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3133_addr_0
    process(ptr_deref_3133_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3133_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3133_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3133_base_resize
    process(arrayidx993_3131) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx993_3131;
      ov := iv(13 downto 0);
      ptr_deref_3133_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3133_gather_scatter
    process(tmp989_3110) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp989_3110;
      ov(63 downto 0) := iv;
      ptr_deref_3133_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3133_root_address_inst
    process(ptr_deref_3133_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3133_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3133_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3571_addr_0
    process(ptr_deref_3571_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3571_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3571_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3571_base_resize
    process(arrayidx1168_3569) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1168_3569;
      ov := iv(13 downto 0);
      ptr_deref_3571_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3571_gather_scatter
    process(type_cast_3573_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3573_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3571_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3571_root_address_inst
    process(ptr_deref_3571_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3571_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3571_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3655_addr_0
    process(ptr_deref_3655_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3655_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3655_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3655_base_resize
    process(arrayidx1211_3652) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1211_3652;
      ov := iv(13 downto 0);
      ptr_deref_3655_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3655_gather_scatter
    process(ptr_deref_3655_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3655_data_0;
      ov(63 downto 0) := iv;
      tmp1212_3656 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3655_root_address_inst
    process(ptr_deref_3655_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3655_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3655_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3679_addr_0
    process(ptr_deref_3679_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3679_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3679_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3679_base_resize
    process(arrayidx1216_3677) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1216_3677;
      ov := iv(13 downto 0);
      ptr_deref_3679_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3679_gather_scatter
    process(tmp1212_3656) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1212_3656;
      ov(63 downto 0) := iv;
      ptr_deref_3679_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3679_root_address_inst
    process(ptr_deref_3679_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3679_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3679_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4097_addr_0
    process(ptr_deref_4097_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4097_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4097_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4097_base_resize
    process(arrayidx1386_4095) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1386_4095;
      ov := iv(13 downto 0);
      ptr_deref_4097_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4097_gather_scatter
    process(type_cast_4099_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_4099_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_4097_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4097_root_address_inst
    process(ptr_deref_4097_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4097_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4097_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4181_addr_0
    process(ptr_deref_4181_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4181_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4181_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4181_base_resize
    process(arrayidx1429_4178) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1429_4178;
      ov := iv(13 downto 0);
      ptr_deref_4181_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4181_gather_scatter
    process(ptr_deref_4181_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4181_data_0;
      ov(63 downto 0) := iv;
      tmp1430_4182 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4181_root_address_inst
    process(ptr_deref_4181_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4181_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4181_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4205_addr_0
    process(ptr_deref_4205_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4205_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4205_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4205_base_resize
    process(arrayidx1434_4203) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1434_4203;
      ov := iv(13 downto 0);
      ptr_deref_4205_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4205_gather_scatter
    process(tmp1430_4182) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1430_4182;
      ov(63 downto 0) := iv;
      ptr_deref_4205_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4205_root_address_inst
    process(ptr_deref_4205_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4205_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4205_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4625_addr_0
    process(ptr_deref_4625_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4625_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4625_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4625_base_resize
    process(arrayidx1606_4623) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1606_4623;
      ov := iv(13 downto 0);
      ptr_deref_4625_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4625_gather_scatter
    process(type_cast_4627_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_4627_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_4625_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4625_root_address_inst
    process(ptr_deref_4625_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4625_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4625_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4709_addr_0
    process(ptr_deref_4709_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4709_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4709_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4709_base_resize
    process(arrayidx1649_4706) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1649_4706;
      ov := iv(13 downto 0);
      ptr_deref_4709_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4709_gather_scatter
    process(ptr_deref_4709_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4709_data_0;
      ov(63 downto 0) := iv;
      tmp1650_4710 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4709_root_address_inst
    process(ptr_deref_4709_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4709_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4709_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4733_addr_0
    process(ptr_deref_4733_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4733_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4733_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4733_base_resize
    process(arrayidx1654_4731) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1654_4731;
      ov := iv(13 downto 0);
      ptr_deref_4733_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4733_gather_scatter
    process(tmp1650_4710) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1650_4710;
      ov(63 downto 0) := iv;
      ptr_deref_4733_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4733_root_address_inst
    process(ptr_deref_4733_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4733_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4733_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_924_addr_0
    process(ptr_deref_924_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_924_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_924_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_924_base_resize
    process(arrayidx_922) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_922;
      ov := iv(13 downto 0);
      ptr_deref_924_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_924_gather_scatter
    process(type_cast_926_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_926_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_924_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_924_root_address_inst
    process(ptr_deref_924_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_924_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_924_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1055_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp133_1054;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1055_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1055_branch_req_0,
          ack0 => if_stmt_1055_branch_ack_0,
          ack1 => if_stmt_1055_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1148_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp166_1147;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1148_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1148_branch_req_0,
          ack0 => if_stmt_1148_branch_ack_0,
          ack1 => if_stmt_1148_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1309_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp239_1308;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1309_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1309_branch_req_0,
          ack0 => if_stmt_1309_branch_ack_0,
          ack1 => if_stmt_1309_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1341_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp250_1340;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1341_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1341_branch_req_0,
          ack0 => if_stmt_1341_branch_ack_0,
          ack1 => if_stmt_1341_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1360_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp257_1359;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1360_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1360_branch_req_0,
          ack0 => if_stmt_1360_branch_ack_0,
          ack1 => if_stmt_1360_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1386_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp267_1385;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1386_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1386_branch_req_0,
          ack0 => if_stmt_1386_branch_ack_0,
          ack1 => if_stmt_1386_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1576_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp346_1575;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1576_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1576_branch_req_0,
          ack0 => if_stmt_1576_branch_ack_0,
          ack1 => if_stmt_1576_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1662_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp380_1661;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1662_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1662_branch_req_0,
          ack0 => if_stmt_1662_branch_ack_0,
          ack1 => if_stmt_1662_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1823_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp455_1822;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1823_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1823_branch_req_0,
          ack0 => if_stmt_1823_branch_ack_0,
          ack1 => if_stmt_1823_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1855_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp466_1854;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1855_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1855_branch_req_0,
          ack0 => if_stmt_1855_branch_ack_0,
          ack1 => if_stmt_1855_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1874_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp473_1873;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1874_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1874_branch_req_0,
          ack0 => if_stmt_1874_branch_ack_0,
          ack1 => if_stmt_1874_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1906_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp484_1905;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1906_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1906_branch_req_0,
          ack0 => if_stmt_1906_branch_ack_0,
          ack1 => if_stmt_1906_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2096_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp563_2095;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2096_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2096_branch_req_0,
          ack0 => if_stmt_2096_branch_ack_0,
          ack1 => if_stmt_2096_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2189_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp598_2188;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2189_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2189_branch_req_0,
          ack0 => if_stmt_2189_branch_ack_0,
          ack1 => if_stmt_2189_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2363_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp677_2362;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2363_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2363_branch_req_0,
          ack0 => if_stmt_2363_branch_ack_0,
          ack1 => if_stmt_2363_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2395_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp688_2394;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2395_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2395_branch_req_0,
          ack0 => if_stmt_2395_branch_ack_0,
          ack1 => if_stmt_2395_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2414_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp695_2413;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2414_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2414_branch_req_0,
          ack0 => if_stmt_2414_branch_ack_0,
          ack1 => if_stmt_2414_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2440_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp705_2439;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2440_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2440_branch_req_0,
          ack0 => if_stmt_2440_branch_ack_0,
          ack1 => if_stmt_2440_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2630_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp784_2629;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2630_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2630_branch_req_0,
          ack0 => if_stmt_2630_branch_ack_0,
          ack1 => if_stmt_2630_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2716_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp818_2715;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2716_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2716_branch_req_0,
          ack0 => if_stmt_2716_branch_ack_0,
          ack1 => if_stmt_2716_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2877_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp893_2876;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2877_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2877_branch_req_0,
          ack0 => if_stmt_2877_branch_ack_0,
          ack1 => if_stmt_2877_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2915_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp905_2914;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2915_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2915_branch_req_0,
          ack0 => if_stmt_2915_branch_ack_0,
          ack1 => if_stmt_2915_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2934_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp912_2933;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2934_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2934_branch_req_0,
          ack0 => if_stmt_2934_branch_ack_0,
          ack1 => if_stmt_2934_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2966_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp923_2965;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2966_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2966_branch_req_0,
          ack0 => if_stmt_2966_branch_ack_0,
          ack1 => if_stmt_2966_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3156_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1002_3155;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3156_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3156_branch_req_0,
          ack0 => if_stmt_3156_branch_ack_0,
          ack1 => if_stmt_3156_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3255_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1038_3254;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3255_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3255_branch_req_0,
          ack0 => if_stmt_3255_branch_ack_0,
          ack1 => if_stmt_3255_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3429_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1117_3428;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3429_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3429_branch_req_0,
          ack0 => if_stmt_3429_branch_ack_0,
          ack1 => if_stmt_3429_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3467_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1129_3466;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3467_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3467_branch_req_0,
          ack0 => if_stmt_3467_branch_ack_0,
          ack1 => if_stmt_3467_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3486_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1136_3485;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3486_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3486_branch_req_0,
          ack0 => if_stmt_3486_branch_ack_0,
          ack1 => if_stmt_3486_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3512_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1146_3511;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3512_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3512_branch_req_0,
          ack0 => if_stmt_3512_branch_ack_0,
          ack1 => if_stmt_3512_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3702_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1225_3701;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3702_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3702_branch_req_0,
          ack0 => if_stmt_3702_branch_ack_0,
          ack1 => if_stmt_3702_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3794_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1260_3793;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3794_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3794_branch_req_0,
          ack0 => if_stmt_3794_branch_ack_0,
          ack1 => if_stmt_3794_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3961_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1336_3960;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3961_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3961_branch_req_0,
          ack0 => if_stmt_3961_branch_ack_0,
          ack1 => if_stmt_3961_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3987_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1346_3986;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3987_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3987_branch_req_0,
          ack0 => if_stmt_3987_branch_ack_0,
          ack1 => if_stmt_3987_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4006_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1353_4005;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4006_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4006_branch_req_0,
          ack0 => if_stmt_4006_branch_ack_0,
          ack1 => if_stmt_4006_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4038_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1364_4037;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4038_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4038_branch_req_0,
          ack0 => if_stmt_4038_branch_ack_0,
          ack1 => if_stmt_4038_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4228_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1443_4227;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4228_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4228_branch_req_0,
          ack0 => if_stmt_4228_branch_ack_0,
          ack1 => if_stmt_4228_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4315_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1477_4314;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4315_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4315_branch_req_0,
          ack0 => if_stmt_4315_branch_ack_0,
          ack1 => if_stmt_4315_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4495_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1557_4494;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4495_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4495_branch_req_0,
          ack0 => if_stmt_4495_branch_ack_0,
          ack1 => if_stmt_4495_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4521_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1567_4520;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4521_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4521_branch_req_0,
          ack0 => if_stmt_4521_branch_ack_0,
          ack1 => if_stmt_4521_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4540_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1574_4539;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4540_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4540_branch_req_0,
          ack0 => if_stmt_4540_branch_ack_0,
          ack1 => if_stmt_4540_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4566_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1584_4565;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4566_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4566_branch_req_0,
          ack0 => if_stmt_4566_branch_ack_0,
          ack1 => if_stmt_4566_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4756_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1663_4755;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4756_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4756_branch_req_0,
          ack0 => if_stmt_4756_branch_ack_0,
          ack1 => if_stmt_4756_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4836_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1696_4835;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4836_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4836_branch_req_0,
          ack0 => if_stmt_4836_branch_ack_0,
          ack1 => if_stmt_4836_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_781_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_780;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_781_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_781_branch_req_0,
          ack0 => if_stmt_781_branch_ack_0,
          ack1 => if_stmt_781_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_813_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp46_812;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_813_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_813_branch_req_0,
          ack0 => if_stmt_813_branch_ack_0,
          ack1 => if_stmt_813_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_832_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp53_831;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_832_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_832_branch_req_0,
          ack0 => if_stmt_832_branch_ack_0,
          ack1 => if_stmt_832_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_864_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp64_863;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_864_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_864_branch_req_0,
          ack0 => if_stmt_864_branch_ack_0,
          ack1 => if_stmt_864_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1066_inst
    process(kx_x1_761) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_761, type_cast_1065_wire_constant, tmp_var);
      add138_1067 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1074_inst
    process(jx_x1_747) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_747, type_cast_1073_wire_constant, tmp_var);
      inc_1075 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1111_inst
    process(inc155_1107, ix_x2_754) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc155_1107, ix_x2_754, tmp_var);
      inc155x_xix_x2_1112 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1587_inst
    process(k176x_x1_1289) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k176x_x1_1289, type_cast_1586_wire_constant, tmp_var);
      add351_1588 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1595_inst
    process(j230x_x1_1276) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j230x_x1_1276, type_cast_1594_wire_constant, tmp_var);
      inc355_1596 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1626_inst
    process(inc369_1622, i184x_x2_1282) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc369_1622, i184x_x2_1282, tmp_var);
      inc369x_xi184x_x2_1627 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2107_inst
    process(k392x_x1_1790) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k392x_x1_1790, type_cast_2106_wire_constant, tmp_var);
      add568_2108 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2115_inst
    process(j446x_x1_1803) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j446x_x1_1803, type_cast_2114_wire_constant, tmp_var);
      inc572_2116 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2152_inst
    process(inc587_2148, i396x_x2_1797) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc587_2148, i396x_x2_1797, tmp_var);
      inc587x_xi396x_x2_2153 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2641_inst
    process(k610x_x1_2331) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k610x_x1_2331, type_cast_2640_wire_constant, tmp_var);
      add789_2642 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2649_inst
    process(j668x_x1_2344) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j668x_x1_2344, type_cast_2648_wire_constant, tmp_var);
      inc793_2650 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2680_inst
    process(inc807_2676, i618x_x2_2338) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc807_2676, i618x_x2_2338, tmp_var);
      inc807x_xi618x_x2_2681 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3167_inst
    process(k830x_x1_2844) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k830x_x1_2844, type_cast_3166_wire_constant, tmp_var);
      add1007_3168 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3175_inst
    process(j884x_x1_2857) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j884x_x1_2857, type_cast_3174_wire_constant, tmp_var);
      inc1011_3176 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3212_inst
    process(inc1026_3208, i834x_x2_2851) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1026_3208, i834x_x2_2851, tmp_var);
      inc1026x_xi834x_x2_3213 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3713_inst
    process(k1050x_x1_3397) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1050x_x1_3397, type_cast_3712_wire_constant, tmp_var);
      add1230_3714 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3721_inst
    process(j1108x_x1_3410) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1108x_x1_3410, type_cast_3720_wire_constant, tmp_var);
      inc1234_3722 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3752_inst
    process(inc1248_3748, i1058x_x2_3404) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1248_3748, i1058x_x2_3404, tmp_var);
      inc1248x_xi1058x_x2_3753 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4239_inst
    process(k1272x_x1_3928) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1272x_x1_3928, type_cast_4238_wire_constant, tmp_var);
      add1448_4240 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4247_inst
    process(j1327x_x1_3941) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1327x_x1_3941, type_cast_4246_wire_constant, tmp_var);
      inc1452_4248 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4284_inst
    process(inc1467_4280, i1276x_x2_3935) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1467_4280, i1276x_x2_3935, tmp_var);
      inc1467x_xi1276x_x2_4285 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4767_inst
    process(k1489x_x1_4463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1489x_x1_4463, type_cast_4766_wire_constant, tmp_var);
      add1668_4768 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4775_inst
    process(j1548x_x1_4476) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1548x_x1_4476, type_cast_4774_wire_constant, tmp_var);
      inc1672_4776 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4806_inst
    process(inc1686_4802, i1497x_x2_4470) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1686_4802, i1497x_x2_4470, tmp_var);
      inc1686x_xi1497x_x2_4807 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1046_inst
    process(conv129_1041) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv129_1041, type_cast_1045_wire_constant, tmp_var);
      add130_1047 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1097_inst
    process(div146_1093, shl_724) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div146_1093, shl_724, tmp_var);
      add149_1098 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1141_inst
    process(div161_1137, shl_724) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div161_1137, shl_724, tmp_var);
      add165_1142 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1332_inst
    process(div246_1328, conv238_1228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div246_1328, conv238_1228, tmp_var);
      add249_1333 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1377_inst
    process(conv263_1373, conv238_1228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv263_1373, conv238_1228, tmp_var);
      add266_1378 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1416_inst
    process(mul284_1412, mul278_1407) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul284_1412, mul278_1407, tmp_var);
      add279_1417 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1421_inst
    process(add279_1417, conv273_1397) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add279_1417, conv273_1397, tmp_var);
      add285_1422 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1479_inst
    process(conv294_1455, mul302_1465) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv294_1455, mul302_1465, tmp_var);
      add303_1480 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1484_inst
    process(add303_1480, mul311_1475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add303_1480, mul311_1475, tmp_var);
      add312_1485 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1499_inst
    process(mul327_1495, mul321_1490) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul327_1495, mul321_1490, tmp_var);
      add322_1500 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1504_inst
    process(add322_1500, conv294_1455) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add322_1500, conv294_1455, tmp_var);
      add328_1505 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1567_inst
    process(conv342_1562) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv342_1562, type_cast_1566_wire_constant, tmp_var);
      add343_1568 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1612_inst
    process(conv359_1608, shl362_1253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv359_1608, shl362_1253, tmp_var);
      add363_1613 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1655_inst
    process(div375_1651, shl362_1253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div375_1651, shl362_1253, tmp_var);
      add379_1656 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1846_inst
    process(div462_1842, conv454_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div462_1842, conv454_1742, tmp_var);
      add465_1847 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1897_inst
    process(div480_1893, conv454_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div480_1893, conv454_1742, tmp_var);
      add483_1898 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1936_inst
    process(mul501_1932, conv490_1917) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul501_1932, conv490_1917, tmp_var);
      add496_1937 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1941_inst
    process(add496_1937, mul495_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add496_1937, mul495_1927, tmp_var);
      add502_1942 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1999_inst
    process(mul528_1995, conv511_1975) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul528_1995, conv511_1975, tmp_var);
      add520_2000 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2004_inst
    process(add520_2000, mul519_1985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add520_2000, mul519_1985, tmp_var);
      add529_2005 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2019_inst
    process(mul544_2015, conv511_1975) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul544_2015, conv511_1975, tmp_var);
      add539_2020 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2024_inst
    process(add539_2020, mul538_2010) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add539_2020, mul538_2010, tmp_var);
      add545_2025 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2087_inst
    process(conv559_2082) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv559_2082, type_cast_2086_wire_constant, tmp_var);
      add560_2088 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2138_inst
    process(div577_2134, shl580_1767) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div577_2134, shl580_1767, tmp_var);
      add581_2139 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2182_inst
    process(div593_2178, shl580_1767) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div593_2178, shl580_1767, tmp_var);
      add597_2183 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2386_inst
    process(div684_2382, conv676_2283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div684_2382, conv676_2283, tmp_var);
      add687_2387 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2431_inst
    process(conv701_2427, conv676_2283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv701_2427, conv676_2283, tmp_var);
      add704_2432 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2470_inst
    process(mul722_2466, conv711_2451) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul722_2466, conv711_2451, tmp_var);
      add717_2471 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2475_inst
    process(add717_2471, mul716_2461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add717_2471, mul716_2461, tmp_var);
      add723_2476 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2533_inst
    process(mul749_2529, conv732_2509) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul749_2529, conv732_2509, tmp_var);
      add741_2534 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2538_inst
    process(add741_2534, mul740_2519) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add741_2534, mul740_2519, tmp_var);
      add750_2539 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2553_inst
    process(mul765_2549, conv732_2509) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul765_2549, conv732_2509, tmp_var);
      add760_2554 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2558_inst
    process(add760_2554, mul759_2544) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add760_2554, mul759_2544, tmp_var);
      add766_2559 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2621_inst
    process(conv780_2616) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv780_2616, type_cast_2620_wire_constant, tmp_var);
      add781_2622 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2666_inst
    process(conv797_2662, shl800_2308) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv797_2662, shl800_2308, tmp_var);
      add801_2667 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2709_inst
    process(div813_2705, shl800_2308) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div813_2705, shl800_2308, tmp_var);
      add817_2710 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2906_inst
    process(div901_2902, conv892_2796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div901_2902, conv892_2796, tmp_var);
      add904_2907 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2957_inst
    process(div919_2953, conv892_2796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div919_2953, conv892_2796, tmp_var);
      add922_2958 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2996_inst
    process(mul940_2992, conv929_2977) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul940_2992, conv929_2977, tmp_var);
      add935_2997 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3001_inst
    process(add935_2997, mul934_2987) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add935_2997, mul934_2987, tmp_var);
      add941_3002 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3059_inst
    process(mul967_3055, conv950_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul967_3055, conv950_3035, tmp_var);
      add959_3060 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3064_inst
    process(add959_3060, mul958_3045) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add959_3060, mul958_3045, tmp_var);
      add968_3065 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3079_inst
    process(mul983_3075, conv950_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul983_3075, conv950_3035, tmp_var);
      add978_3080 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3084_inst
    process(add978_3080, mul977_3070) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add978_3080, mul977_3070, tmp_var);
      add984_3085 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3147_inst
    process(conv998_3142) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv998_3142, type_cast_3146_wire_constant, tmp_var);
      add999_3148 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3198_inst
    process(div1016_3194, shl1019_2821) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1016_3194, shl1019_2821, tmp_var);
      add1020_3199 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3248_inst
    process(div1033_3244, shl1019_2821) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1033_3244, shl1019_2821, tmp_var);
      add1037_3249 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3458_inst
    process(div1125_3454, conv1116_3349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1125_3454, conv1116_3349, tmp_var);
      add1128_3459 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3503_inst
    process(conv1142_3499, conv1116_3349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1142_3499, conv1116_3349, tmp_var);
      add1145_3504 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3542_inst
    process(mul1163_3538, conv1152_3523) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1163_3538, conv1152_3523, tmp_var);
      add1158_3543 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3547_inst
    process(add1158_3543, mul1157_3533) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1158_3543, mul1157_3533, tmp_var);
      add1164_3548 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3605_inst
    process(mul1190_3601, conv1173_3581) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1190_3601, conv1173_3581, tmp_var);
      add1182_3606 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3610_inst
    process(add1182_3606, mul1181_3591) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1182_3606, mul1181_3591, tmp_var);
      add1191_3611 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3625_inst
    process(mul1206_3621, conv1173_3581) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1206_3621, conv1173_3581, tmp_var);
      add1201_3626 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3630_inst
    process(add1201_3626, mul1200_3616) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1201_3626, mul1200_3616, tmp_var);
      add1207_3631 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3693_inst
    process(conv1221_3688) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1221_3688, type_cast_3692_wire_constant, tmp_var);
      add1222_3694 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3738_inst
    process(conv1238_3734, shl1241_3374) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1238_3734, shl1241_3374, tmp_var);
      add1242_3739 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3787_inst
    process(div1255_3783, shl1241_3374) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1255_3783, shl1241_3374, tmp_var);
      add1259_3788 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3978_inst
    process(conv1342_3974, conv1335_3880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1342_3974, conv1335_3880, tmp_var);
      add1345_3979 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4029_inst
    process(div1360_4025, conv1335_3880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1360_4025, conv1335_3880, tmp_var);
      add1363_4030 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4068_inst
    process(mul1381_4064, conv1370_4049) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1381_4064, conv1370_4049, tmp_var);
      add1376_4069 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4073_inst
    process(add1376_4069, mul1375_4059) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1376_4069, mul1375_4059, tmp_var);
      add1382_4074 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4131_inst
    process(mul1408_4127, conv1391_4107) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1408_4127, conv1391_4107, tmp_var);
      add1400_4132 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4136_inst
    process(add1400_4132, mul1399_4117) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1400_4132, mul1399_4117, tmp_var);
      add1409_4137 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4151_inst
    process(mul1424_4147, conv1391_4107) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1424_4147, conv1391_4107, tmp_var);
      add1419_4152 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4156_inst
    process(add1419_4152, mul1418_4142) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1419_4152, mul1418_4142, tmp_var);
      add1425_4157 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4219_inst
    process(conv1439_4214) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1439_4214, type_cast_4218_wire_constant, tmp_var);
      add1440_4220 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4270_inst
    process(div1457_4266, shl1460_3905) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1457_4266, shl1460_3905, tmp_var);
      add1461_4271 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4308_inst
    process(conv1472_4304, shl1460_3905) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1472_4304, shl1460_3905, tmp_var);
      add1476_4309 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4512_inst
    process(conv1563_4508, conv1556_4415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1563_4508, conv1556_4415, tmp_var);
      add1566_4513 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4557_inst
    process(conv1580_4553, conv1556_4415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1580_4553, conv1556_4415, tmp_var);
      add1583_4558 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4596_inst
    process(mul1601_4592, conv1590_4577) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1601_4592, conv1590_4577, tmp_var);
      add1596_4597 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4601_inst
    process(add1596_4597, mul1595_4587) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1596_4597, mul1595_4587, tmp_var);
      add1602_4602 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4659_inst
    process(mul1628_4655, conv1611_4635) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1628_4655, conv1611_4635, tmp_var);
      add1620_4660 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4664_inst
    process(add1620_4660, mul1619_4645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1620_4660, mul1619_4645, tmp_var);
      add1629_4665 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4679_inst
    process(mul1644_4675, conv1611_4635) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1644_4675, conv1611_4635, tmp_var);
      add1639_4680 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4684_inst
    process(add1639_4680, mul1638_4670) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1639_4680, mul1638_4670, tmp_var);
      add1645_4685 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4747_inst
    process(conv1659_4742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1659_4742, type_cast_4746_wire_constant, tmp_var);
      add1660_4748 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4792_inst
    process(conv1676_4788, shl1679_4440) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1676_4788, shl1679_4440, tmp_var);
      add1680_4793 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4829_inst
    process(conv1691_4825, shl1679_4440) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1691_4825, shl1679_4440, tmp_var);
      add1695_4830 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_804_inst
    process(div_800, conv38_698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div_800, conv38_698, tmp_var);
      add_805 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_855_inst
    process(div60_851, conv38_698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div60_851, conv38_698, tmp_var);
      add63_856 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_894_inst
    process(mul79_890, mul73_885) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul79_890, mul73_885, tmp_var);
      add74_895 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_899_inst
    process(add74_895, conv68_875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_895, conv68_875, tmp_var);
      add80_900 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_958_inst
    process(conv84_934, mul91_944) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv84_934, mul91_944, tmp_var);
      add92_959 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_963_inst
    process(add92_959, mul100_954) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add92_959, mul100_954, tmp_var);
      add101_964 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_978_inst
    process(mul116_974, mul110_969) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul116_974, mul110_969, tmp_var);
      add111_979 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_983_inst
    process(add111_979, conv84_934) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add111_979, conv84_934, tmp_var);
      add117_984 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1016_inst
    process(type_cast_1012_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1012_wire, type_cast_1015_wire_constant, tmp_var);
      ASHR_i32_i32_1016_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1245_inst
    process(type_cast_1241_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1241_wire, type_cast_1244_wire_constant, tmp_var);
      ASHR_i32_i32_1245_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1271_inst
    process(type_cast_1267_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1267_wire, type_cast_1270_wire_constant, tmp_var);
      ASHR_i32_i32_1271_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1429_inst
    process(type_cast_1425_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1425_wire, type_cast_1428_wire_constant, tmp_var);
      ASHR_i32_i32_1429_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1512_inst
    process(type_cast_1508_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1508_wire, type_cast_1511_wire_constant, tmp_var);
      ASHR_i32_i32_1512_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1537_inst
    process(type_cast_1533_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1533_wire, type_cast_1536_wire_constant, tmp_var);
      ASHR_i32_i32_1537_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1759_inst
    process(type_cast_1755_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1755_wire, type_cast_1758_wire_constant, tmp_var);
      ASHR_i32_i32_1759_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1785_inst
    process(type_cast_1781_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1781_wire, type_cast_1784_wire_constant, tmp_var);
      ASHR_i32_i32_1785_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1949_inst
    process(type_cast_1945_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1945_wire, type_cast_1948_wire_constant, tmp_var);
      ASHR_i32_i32_1949_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2032_inst
    process(type_cast_2028_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2028_wire, type_cast_2031_wire_constant, tmp_var);
      ASHR_i32_i32_2032_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2057_inst
    process(type_cast_2053_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2053_wire, type_cast_2056_wire_constant, tmp_var);
      ASHR_i32_i32_2057_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2300_inst
    process(type_cast_2296_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2296_wire, type_cast_2299_wire_constant, tmp_var);
      ASHR_i32_i32_2300_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2326_inst
    process(type_cast_2322_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2322_wire, type_cast_2325_wire_constant, tmp_var);
      ASHR_i32_i32_2326_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2483_inst
    process(type_cast_2479_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2479_wire, type_cast_2482_wire_constant, tmp_var);
      ASHR_i32_i32_2483_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2566_inst
    process(type_cast_2562_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2562_wire, type_cast_2565_wire_constant, tmp_var);
      ASHR_i32_i32_2566_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2591_inst
    process(type_cast_2587_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2587_wire, type_cast_2590_wire_constant, tmp_var);
      ASHR_i32_i32_2591_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2813_inst
    process(type_cast_2809_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2809_wire, type_cast_2812_wire_constant, tmp_var);
      ASHR_i32_i32_2813_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2839_inst
    process(type_cast_2835_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2835_wire, type_cast_2838_wire_constant, tmp_var);
      ASHR_i32_i32_2839_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3009_inst
    process(type_cast_3005_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3005_wire, type_cast_3008_wire_constant, tmp_var);
      ASHR_i32_i32_3009_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3092_inst
    process(type_cast_3088_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3088_wire, type_cast_3091_wire_constant, tmp_var);
      ASHR_i32_i32_3092_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3117_inst
    process(type_cast_3113_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3113_wire, type_cast_3116_wire_constant, tmp_var);
      ASHR_i32_i32_3117_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3366_inst
    process(type_cast_3362_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3362_wire, type_cast_3365_wire_constant, tmp_var);
      ASHR_i32_i32_3366_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3392_inst
    process(type_cast_3388_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3388_wire, type_cast_3391_wire_constant, tmp_var);
      ASHR_i32_i32_3392_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3555_inst
    process(type_cast_3551_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3551_wire, type_cast_3554_wire_constant, tmp_var);
      ASHR_i32_i32_3555_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3638_inst
    process(type_cast_3634_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3634_wire, type_cast_3637_wire_constant, tmp_var);
      ASHR_i32_i32_3638_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3663_inst
    process(type_cast_3659_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3659_wire, type_cast_3662_wire_constant, tmp_var);
      ASHR_i32_i32_3663_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3897_inst
    process(type_cast_3893_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3893_wire, type_cast_3896_wire_constant, tmp_var);
      ASHR_i32_i32_3897_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3923_inst
    process(type_cast_3919_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3919_wire, type_cast_3922_wire_constant, tmp_var);
      ASHR_i32_i32_3923_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4081_inst
    process(type_cast_4077_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4077_wire, type_cast_4080_wire_constant, tmp_var);
      ASHR_i32_i32_4081_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4164_inst
    process(type_cast_4160_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4160_wire, type_cast_4163_wire_constant, tmp_var);
      ASHR_i32_i32_4164_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4189_inst
    process(type_cast_4185_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4185_wire, type_cast_4188_wire_constant, tmp_var);
      ASHR_i32_i32_4189_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4432_inst
    process(type_cast_4428_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4428_wire, type_cast_4431_wire_constant, tmp_var);
      ASHR_i32_i32_4432_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4458_inst
    process(type_cast_4454_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4454_wire, type_cast_4457_wire_constant, tmp_var);
      ASHR_i32_i32_4458_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4609_inst
    process(type_cast_4605_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4605_wire, type_cast_4608_wire_constant, tmp_var);
      ASHR_i32_i32_4609_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4692_inst
    process(type_cast_4688_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4688_wire, type_cast_4691_wire_constant, tmp_var);
      ASHR_i32_i32_4692_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4717_inst
    process(type_cast_4713_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4713_wire, type_cast_4716_wire_constant, tmp_var);
      ASHR_i32_i32_4717_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_716_inst
    process(type_cast_712_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_712_wire, type_cast_715_wire_constant, tmp_var);
      ASHR_i32_i32_716_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_742_inst
    process(type_cast_738_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_738_wire, type_cast_741_wire_constant, tmp_var);
      ASHR_i32_i32_742_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_907_inst
    process(type_cast_903_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_903_wire, type_cast_906_wire_constant, tmp_var);
      ASHR_i32_i32_907_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_991_inst
    process(type_cast_987_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_987_wire, type_cast_990_wire_constant, tmp_var);
      ASHR_i32_i32_991_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1102_inst
    process(conv143_1080, add149_1098) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv143_1080, add149_1098, tmp_var);
      cmp150_1103 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1146_inst
    process(conv158_1124, add165_1142) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv158_1124, add165_1142, tmp_var);
      cmp166_1147 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1617_inst
    process(conv357_1601, add363_1613) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv357_1601, add363_1613, tmp_var);
      cmp364_1618 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1660_inst
    process(conv372_1638, add379_1656) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv372_1638, add379_1656, tmp_var);
      cmp380_1661 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2143_inst
    process(conv574_2121, add581_2139) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv574_2121, add581_2139, tmp_var);
      cmp582_2144 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2187_inst
    process(conv590_2165, add597_2183) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv590_2165, add597_2183, tmp_var);
      cmp598_2188 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2671_inst
    process(conv795_2655, add801_2667) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv795_2655, add801_2667, tmp_var);
      cmp802_2672 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2714_inst
    process(conv810_2692, add817_2710) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv810_2692, add817_2710, tmp_var);
      cmp818_2715 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3203_inst
    process(conv1013_3181, add1020_3199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1013_3181, add1020_3199, tmp_var);
      cmp1021_3204 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3253_inst
    process(conv1029_3225, add1037_3249) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1029_3225, add1037_3249, tmp_var);
      cmp1038_3254 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3743_inst
    process(conv1236_3727, add1242_3739) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1236_3727, add1242_3739, tmp_var);
      cmp1243_3744 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3792_inst
    process(conv1251_3764, add1259_3788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1251_3764, add1259_3788, tmp_var);
      cmp1260_3793 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4275_inst
    process(conv1454_4253, add1461_4271) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1454_4253, add1461_4271, tmp_var);
      cmp1462_4276 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4313_inst
    process(conv1470_4297, add1476_4309) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1470_4297, add1476_4309, tmp_var);
      cmp1477_4314 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4797_inst
    process(conv1674_4781, add1680_4793) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1674_4781, add1680_4793, tmp_var);
      cmp1681_4798 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4834_inst
    process(conv1689_4818, add1695_4830) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1689_4818, add1695_4830, tmp_var);
      cmp1696_4835 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1194_inst
    process(conv180_1189) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv180_1189, type_cast_1193_wire_constant, tmp_var);
      div181_1195 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1708_inst
    process(conv398_1703) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv398_1703, type_cast_1707_wire_constant, tmp_var);
      div399_1709 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2239_inst
    process(conv614_2234) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv614_2234, type_cast_2238_wire_constant, tmp_var);
      div615_2240 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2249_inst
    process(conv620_2244) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv620_2244, type_cast_2248_wire_constant, tmp_var);
      div621_2250 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2762_inst
    process(conv836_2757) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv836_2757, type_cast_2761_wire_constant, tmp_var);
      div837_2763 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3305_inst
    process(conv1054_3300) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1054_3300, type_cast_3304_wire_constant, tmp_var);
      div1055_3306 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3315_inst
    process(conv1060_3310) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1060_3310, type_cast_3314_wire_constant, tmp_var);
      div1061_3316 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3840_inst
    process(conv1278_3835) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1278_3835, type_cast_3839_wire_constant, tmp_var);
      div1279_3841 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4365_inst
    process(conv1493_4360) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1493_4360, type_cast_4364_wire_constant, tmp_var);
      div1494_4366 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4381_inst
    process(mul1500_4376) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1500_4376, type_cast_4380_wire_constant, tmp_var);
      div1501_4382 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1092_inst
    process(conv145_1087) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv145_1087, type_cast_1091_wire_constant, tmp_var);
      div146_1093 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1136_inst
    process(conv160_1131) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv160_1131, type_cast_1135_wire_constant, tmp_var);
      div161_1137 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1327_inst
    process(conv245_1322) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv245_1322, type_cast_1326_wire_constant, tmp_var);
      div246_1328 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1650_inst
    process(conv374_1645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv374_1645, type_cast_1649_wire_constant, tmp_var);
      div375_1651 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1841_inst
    process(conv461_1836) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv461_1836, type_cast_1840_wire_constant, tmp_var);
      div462_1842 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1892_inst
    process(conv479_1887) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv479_1887, type_cast_1891_wire_constant, tmp_var);
      div480_1893 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2133_inst
    process(conv576_2128) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv576_2128, type_cast_2132_wire_constant, tmp_var);
      div577_2134 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2177_inst
    process(conv592_2172) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv592_2172, type_cast_2176_wire_constant, tmp_var);
      div593_2178 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2381_inst
    process(conv683_2376) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv683_2376, type_cast_2380_wire_constant, tmp_var);
      div684_2382 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2704_inst
    process(conv812_2699) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv812_2699, type_cast_2703_wire_constant, tmp_var);
      div813_2705 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2901_inst
    process(mul900_2896) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul900_2896, type_cast_2900_wire_constant, tmp_var);
      div901_2902 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2952_inst
    process(conv918_2947) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv918_2947, type_cast_2951_wire_constant, tmp_var);
      div919_2953 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3193_inst
    process(conv1015_3188) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1015_3188, type_cast_3192_wire_constant, tmp_var);
      div1016_3194 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3243_inst
    process(mul1032_3238) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1032_3238, type_cast_3242_wire_constant, tmp_var);
      div1033_3244 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3453_inst
    process(mul1124_3448) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1124_3448, type_cast_3452_wire_constant, tmp_var);
      div1125_3454 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3782_inst
    process(mul1254_3777) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1254_3777, type_cast_3781_wire_constant, tmp_var);
      div1255_3783 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_4024_inst
    process(conv1359_4019) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1359_4019, type_cast_4023_wire_constant, tmp_var);
      div1360_4025 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_4265_inst
    process(conv1456_4260) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1456_4260, type_cast_4264_wire_constant, tmp_var);
      div1457_4266 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_799_inst
    process(conv43_794) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv43_794, type_cast_798_wire_constant, tmp_var);
      div_800 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_850_inst
    process(conv59_845) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv59_845, type_cast_849_wire_constant, tmp_var);
      div60_851 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3846_inst
    process(div1279_3841) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(div1279_3841, type_cast_3845_wire_constant, tmp_var);
      mul1280_3847 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_4375_inst
    process(conv1499_4370) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1499_4370, type_cast_4374_wire_constant, tmp_var);
      mul1500_4376 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1223_inst
    process(conv226_1219, conv224_1215) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv226_1219, conv224_1215, tmp_var);
      mul227_1224 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1263_inst
    process(mul219_1259, conv216_1211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul219_1259, conv216_1211, tmp_var);
      sext1707_1264 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1406_inst
    process(conv277_1402, conv275_1232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv277_1402, conv275_1232, tmp_var);
      mul278_1407 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1411_inst
    process(conv236_1301, conv281_1247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv236_1301, conv281_1247, tmp_var);
      mul284_1412 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1464_inst
    process(sub301_1460, conv216_1211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub301_1460, conv216_1211, tmp_var);
      mul302_1465 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1474_inst
    process(sub310_1470, conv305_1273) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub310_1470, conv305_1273, tmp_var);
      mul311_1475 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1489_inst
    process(conv254_1352, conv275_1232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv254_1352, conv275_1232, tmp_var);
      mul321_1490 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1494_inst
    process(conv236_1301, conv281_1247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv236_1301, conv281_1247, tmp_var);
      mul327_1495 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1737_inst
    process(conv442_1733, conv440_1729) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv442_1733, conv440_1729, tmp_var);
      mul443_1738 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1777_inst
    process(mul435_1773, conv359x_xlcssa_1695) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul435_1773, conv359x_xlcssa_1695, tmp_var);
      sext1708_1778 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1926_inst
    process(conv494_1922, conv492_1746) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv494_1922, conv492_1746, tmp_var);
      mul495_1927 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1931_inst
    process(conv452_1815, conv498_1761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv452_1815, conv498_1761, tmp_var);
      mul501_1932 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1984_inst
    process(sub518_1980, conv432_1725) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub518_1980, conv432_1725, tmp_var);
      mul519_1985 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1994_inst
    process(sub527_1990, conv522_1787) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub527_1990, conv522_1787, tmp_var);
      mul528_1995 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2009_inst
    process(conv470_1866, conv492_1746) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv470_1866, conv492_1746, tmp_var);
      mul538_2010 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2014_inst
    process(conv452_1815, conv498_1761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv452_1815, conv498_1761, tmp_var);
      mul544_2015 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2278_inst
    process(conv664_2274, conv662_2270) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv664_2274, conv662_2270, tmp_var);
      mul665_2279 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2318_inst
    process(mul657_2314, conv576x_xlcssa_2222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul657_2314, conv576x_xlcssa_2222, tmp_var);
      sext1709_2319 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2460_inst
    process(conv715_2456, conv713_2287) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv715_2456, conv713_2287, tmp_var);
      mul716_2461 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2465_inst
    process(conv674_2355, conv719_2302) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv674_2355, conv719_2302, tmp_var);
      mul722_2466 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2518_inst
    process(sub739_2514, conv654_2266) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub739_2514, conv654_2266, tmp_var);
      mul740_2519 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2528_inst
    process(sub748_2524, conv743_2328) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub748_2524, conv743_2328, tmp_var);
      mul749_2529 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2543_inst
    process(conv692_2406, conv713_2287) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv692_2406, conv713_2287, tmp_var);
      mul759_2544 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2548_inst
    process(conv674_2355, conv719_2302) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv674_2355, conv719_2302, tmp_var);
      mul765_2549 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2791_inst
    process(conv880_2787, conv878_2783) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv880_2787, conv878_2783, tmp_var);
      mul881_2792 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2831_inst
    process(mul873_2827, conv797x_xlcssa_2749) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul873_2827, conv797x_xlcssa_2749, tmp_var);
      sext1710_2832 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2895_inst
    process(conv899_2890) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv899_2890, type_cast_2894_wire_constant, tmp_var);
      mul900_2896 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2986_inst
    process(conv933_2982, conv931_2800) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv933_2982, conv931_2800, tmp_var);
      mul934_2987 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2991_inst
    process(conv890_2869, conv937_2815) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv890_2869, conv937_2815, tmp_var);
      mul940_2992 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3044_inst
    process(sub957_3040, conv870_2779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub957_3040, conv870_2779, tmp_var);
      mul958_3045 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3054_inst
    process(sub966_3050, conv961_2841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub966_3050, conv961_2841, tmp_var);
      mul967_3055 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3069_inst
    process(conv909_2926, conv931_2800) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv909_2926, conv931_2800, tmp_var);
      mul977_3070 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3074_inst
    process(conv890_2869, conv937_2815) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv890_2869, conv937_2815, tmp_var);
      mul983_3075 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3237_inst
    process(conv1031_3232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1031_3232, type_cast_3236_wire_constant, tmp_var);
      mul1032_3238 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3344_inst
    process(conv1104_3340, conv1102_3336) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1104_3340, conv1102_3336, tmp_var);
      mul1105_3345 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3384_inst
    process(mul1097_3380, conv1015x_xlcssa_3288) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1097_3380, conv1015x_xlcssa_3288, tmp_var);
      sext1711_3385 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3447_inst
    process(conv1123_3442) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1123_3442, type_cast_3446_wire_constant, tmp_var);
      mul1124_3448 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3532_inst
    process(conv1156_3528, conv1154_3353) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1156_3528, conv1154_3353, tmp_var);
      mul1157_3533 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3537_inst
    process(conv1114_3421, conv1160_3368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1114_3421, conv1160_3368, tmp_var);
      mul1163_3538 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3590_inst
    process(sub1180_3586, conv1094_3332) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1180_3586, conv1094_3332, tmp_var);
      mul1181_3591 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3600_inst
    process(sub1189_3596, conv1184_3394) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1189_3596, conv1184_3394, tmp_var);
      mul1190_3601 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3615_inst
    process(conv1133_3478, conv1154_3353) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1133_3478, conv1154_3353, tmp_var);
      mul1200_3616 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3620_inst
    process(conv1114_3421, conv1160_3368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1114_3421, conv1160_3368, tmp_var);
      mul1206_3621 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3776_inst
    process(conv1253_3771) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1253_3771, type_cast_3775_wire_constant, tmp_var);
      mul1254_3777 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3875_inst
    process(conv1323_3871, conv1321_3867) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1323_3871, conv1321_3867, tmp_var);
      mul1324_3876 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3915_inst
    process(mul1316_3911, conv1238x_xlcssa_3827) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1316_3911, conv1238x_xlcssa_3827, tmp_var);
      sext1712_3916 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4058_inst
    process(conv1374_4054, conv1372_3884) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1374_4054, conv1372_3884, tmp_var);
      mul1375_4059 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4063_inst
    process(conv1333_3953, conv1378_3899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1333_3953, conv1378_3899, tmp_var);
      mul1381_4064 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4116_inst
    process(sub1398_4112, conv1313_3863) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1398_4112, conv1313_3863, tmp_var);
      mul1399_4117 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4126_inst
    process(sub1407_4122, conv1402_3925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1407_4122, conv1402_3925, tmp_var);
      mul1408_4127 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4141_inst
    process(conv1350_3998, conv1372_3884) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1350_3998, conv1372_3884, tmp_var);
      mul1418_4142 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4146_inst
    process(conv1333_3953, conv1378_3899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1333_3953, conv1378_3899, tmp_var);
      mul1424_4147 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4410_inst
    process(conv1544_4406, conv1542_4402) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1544_4406, conv1542_4402, tmp_var);
      mul1545_4411 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4450_inst
    process(mul1537_4446, conv1456x_xlcssa_4348) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1537_4446, conv1456x_xlcssa_4348, tmp_var);
      sext1713_4451 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4586_inst
    process(conv1594_4582, conv1592_4419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1594_4582, conv1592_4419, tmp_var);
      mul1595_4587 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4591_inst
    process(conv1554_4487, conv1598_4434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1554_4487, conv1598_4434, tmp_var);
      mul1601_4592 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4644_inst
    process(sub1618_4640, conv1534_4398) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1618_4640, conv1534_4398, tmp_var);
      mul1619_4645 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4654_inst
    process(sub1627_4650, conv1622_4460) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1627_4650, conv1622_4460, tmp_var);
      mul1628_4655 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4669_inst
    process(conv1571_4532, conv1592_4419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1571_4532, conv1592_4419, tmp_var);
      mul1638_4670 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4674_inst
    process(conv1554_4487, conv1598_4434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1554_4487, conv1598_4434, tmp_var);
      mul1644_4675 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_693_inst
    process(conv29_689, conv27_685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv29_689, conv27_685, tmp_var);
      mul30_694 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_734_inst
    process(mul_730, conv23_681) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_730, conv23_681, tmp_var);
      sext_735 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_884_inst
    process(conv72_880, conv70_702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv72_880, conv70_702, tmp_var);
      mul73_885 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_889_inst
    process(conv36_773, conv76_718) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv36_773, conv76_718, tmp_var);
      mul79_890 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_943_inst
    process(sub_939, conv21_677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_939, conv21_677, tmp_var);
      mul91_944 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_953_inst
    process(sub99_949, conv94_744) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub99_949, conv94_744, tmp_var);
      mul100_954 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_968_inst
    process(conv50_824, conv70_702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv50_824, conv70_702, tmp_var);
      mul110_969 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_973_inst
    process(conv36_773, conv76_718) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv36_773, conv76_718, tmp_var);
      mul116_974 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1237_inst
    process(mul227_1224) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul227_1224, type_cast_1236_wire_constant, tmp_var);
      sext1747_1238 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1252_inst
    process(conv238_1228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv238_1228, type_cast_1251_wire_constant, tmp_var);
      shl362_1253 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1258_inst
    process(conv145x_xlcssa_1177) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv145x_xlcssa_1177, type_cast_1257_wire_constant, tmp_var);
      mul219_1259 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1751_inst
    process(mul443_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul443_1738, type_cast_1750_wire_constant, tmp_var);
      sext1748_1752 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1766_inst
    process(conv454_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv454_1742, type_cast_1765_wire_constant, tmp_var);
      shl580_1767 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1772_inst
    process(conv432_1725) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv432_1725, type_cast_1771_wire_constant, tmp_var);
      mul435_1773 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2292_inst
    process(mul665_2279) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul665_2279, type_cast_2291_wire_constant, tmp_var);
      sext1749_2293 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2307_inst
    process(conv676_2283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv676_2283, type_cast_2306_wire_constant, tmp_var);
      shl800_2308 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2313_inst
    process(conv654_2266) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv654_2266, type_cast_2312_wire_constant, tmp_var);
      mul657_2314 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2805_inst
    process(mul881_2792) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul881_2792, type_cast_2804_wire_constant, tmp_var);
      sext1750_2806 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2820_inst
    process(conv892_2796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv892_2796, type_cast_2819_wire_constant, tmp_var);
      shl1019_2821 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2826_inst
    process(conv870_2779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv870_2779, type_cast_2825_wire_constant, tmp_var);
      mul873_2827 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3358_inst
    process(mul1105_3345) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1105_3345, type_cast_3357_wire_constant, tmp_var);
      sext1751_3359 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3373_inst
    process(conv1116_3349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1116_3349, type_cast_3372_wire_constant, tmp_var);
      shl1241_3374 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3379_inst
    process(conv1094_3332) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1094_3332, type_cast_3378_wire_constant, tmp_var);
      mul1097_3380 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3889_inst
    process(mul1324_3876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1324_3876, type_cast_3888_wire_constant, tmp_var);
      sext1752_3890 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3904_inst
    process(conv1335_3880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1335_3880, type_cast_3903_wire_constant, tmp_var);
      shl1460_3905 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3910_inst
    process(conv1313_3863) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1313_3863, type_cast_3909_wire_constant, tmp_var);
      mul1316_3911 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4424_inst
    process(mul1545_4411) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1545_4411, type_cast_4423_wire_constant, tmp_var);
      sext1753_4425 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4439_inst
    process(conv1556_4415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1556_4415, type_cast_4438_wire_constant, tmp_var);
      shl1679_4440 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4445_inst
    process(conv1534_4398) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1534_4398, type_cast_4444_wire_constant, tmp_var);
      mul1537_4446 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_707_inst
    process(mul30_694) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul30_694, type_cast_706_wire_constant, tmp_var);
      sext1746_708 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_723_inst
    process(conv38_698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv38_698, type_cast_722_wire_constant, tmp_var);
      shl_724 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_729_inst
    process(conv21_677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv21_677, type_cast_728_wire_constant, tmp_var);
      mul_730 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1053_inst
    process(type_cast_1050_wire, type_cast_1052_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1050_wire, type_cast_1052_wire, tmp_var);
      cmp133_1054 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1307_inst
    process(type_cast_1304_wire, type_cast_1306_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1304_wire, type_cast_1306_wire, tmp_var);
      cmp239_1308 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1339_inst
    process(type_cast_1336_wire, type_cast_1338_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1336_wire, type_cast_1338_wire, tmp_var);
      cmp250_1340 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1358_inst
    process(type_cast_1355_wire, type_cast_1357_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1355_wire, type_cast_1357_wire, tmp_var);
      cmp257_1359 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1384_inst
    process(type_cast_1381_wire, type_cast_1383_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1381_wire, type_cast_1383_wire, tmp_var);
      cmp267_1385 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1574_inst
    process(type_cast_1571_wire, type_cast_1573_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1571_wire, type_cast_1573_wire, tmp_var);
      cmp346_1575 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1821_inst
    process(type_cast_1818_wire, type_cast_1820_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1818_wire, type_cast_1820_wire, tmp_var);
      cmp455_1822 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1853_inst
    process(type_cast_1850_wire, type_cast_1852_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1850_wire, type_cast_1852_wire, tmp_var);
      cmp466_1854 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1872_inst
    process(type_cast_1869_wire, type_cast_1871_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1869_wire, type_cast_1871_wire, tmp_var);
      cmp473_1873 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1904_inst
    process(type_cast_1901_wire, type_cast_1903_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1901_wire, type_cast_1903_wire, tmp_var);
      cmp484_1905 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2094_inst
    process(type_cast_2091_wire, type_cast_2093_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2091_wire, type_cast_2093_wire, tmp_var);
      cmp563_2095 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2361_inst
    process(type_cast_2358_wire, type_cast_2360_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2358_wire, type_cast_2360_wire, tmp_var);
      cmp677_2362 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2393_inst
    process(type_cast_2390_wire, type_cast_2392_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2390_wire, type_cast_2392_wire, tmp_var);
      cmp688_2394 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2412_inst
    process(type_cast_2409_wire, type_cast_2411_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2409_wire, type_cast_2411_wire, tmp_var);
      cmp695_2413 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2438_inst
    process(type_cast_2435_wire, type_cast_2437_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2435_wire, type_cast_2437_wire, tmp_var);
      cmp705_2439 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2628_inst
    process(type_cast_2625_wire, type_cast_2627_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2625_wire, type_cast_2627_wire, tmp_var);
      cmp784_2629 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2875_inst
    process(type_cast_2872_wire, type_cast_2874_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2872_wire, type_cast_2874_wire, tmp_var);
      cmp893_2876 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2913_inst
    process(type_cast_2910_wire, type_cast_2912_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2910_wire, type_cast_2912_wire, tmp_var);
      cmp905_2914 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2932_inst
    process(type_cast_2929_wire, type_cast_2931_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2929_wire, type_cast_2931_wire, tmp_var);
      cmp912_2933 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2964_inst
    process(type_cast_2961_wire, type_cast_2963_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2961_wire, type_cast_2963_wire, tmp_var);
      cmp923_2965 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3154_inst
    process(type_cast_3151_wire, type_cast_3153_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3151_wire, type_cast_3153_wire, tmp_var);
      cmp1002_3155 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3427_inst
    process(type_cast_3424_wire, type_cast_3426_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3424_wire, type_cast_3426_wire, tmp_var);
      cmp1117_3428 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3465_inst
    process(type_cast_3462_wire, type_cast_3464_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3462_wire, type_cast_3464_wire, tmp_var);
      cmp1129_3466 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3484_inst
    process(type_cast_3481_wire, type_cast_3483_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3481_wire, type_cast_3483_wire, tmp_var);
      cmp1136_3485 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3510_inst
    process(type_cast_3507_wire, type_cast_3509_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3507_wire, type_cast_3509_wire, tmp_var);
      cmp1146_3511 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3700_inst
    process(type_cast_3697_wire, type_cast_3699_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3697_wire, type_cast_3699_wire, tmp_var);
      cmp1225_3701 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3959_inst
    process(type_cast_3956_wire, type_cast_3958_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3956_wire, type_cast_3958_wire, tmp_var);
      cmp1336_3960 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3985_inst
    process(type_cast_3982_wire, type_cast_3984_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3982_wire, type_cast_3984_wire, tmp_var);
      cmp1346_3986 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4004_inst
    process(type_cast_4001_wire, type_cast_4003_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4001_wire, type_cast_4003_wire, tmp_var);
      cmp1353_4005 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4036_inst
    process(type_cast_4033_wire, type_cast_4035_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4033_wire, type_cast_4035_wire, tmp_var);
      cmp1364_4037 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4226_inst
    process(type_cast_4223_wire, type_cast_4225_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4223_wire, type_cast_4225_wire, tmp_var);
      cmp1443_4227 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4493_inst
    process(type_cast_4490_wire, type_cast_4492_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4490_wire, type_cast_4492_wire, tmp_var);
      cmp1557_4494 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4519_inst
    process(type_cast_4516_wire, type_cast_4518_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4516_wire, type_cast_4518_wire, tmp_var);
      cmp1567_4520 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4538_inst
    process(type_cast_4535_wire, type_cast_4537_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4535_wire, type_cast_4537_wire, tmp_var);
      cmp1574_4539 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4564_inst
    process(type_cast_4561_wire, type_cast_4563_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4561_wire, type_cast_4563_wire, tmp_var);
      cmp1584_4565 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4754_inst
    process(type_cast_4751_wire, type_cast_4753_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4751_wire, type_cast_4753_wire, tmp_var);
      cmp1663_4755 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_779_inst
    process(type_cast_776_wire, type_cast_778_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_776_wire, type_cast_778_wire, tmp_var);
      cmp_780 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_811_inst
    process(type_cast_808_wire, type_cast_810_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_808_wire, type_cast_810_wire, tmp_var);
      cmp46_812 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_830_inst
    process(type_cast_827_wire, type_cast_829_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_827_wire, type_cast_829_wire, tmp_var);
      cmp53_831 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_862_inst
    process(type_cast_859_wire, type_cast_861_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_859_wire, type_cast_861_wire, tmp_var);
      cmp64_863 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1459_inst
    process(conv254_1352, conv238_1228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv254_1352, conv238_1228, tmp_var);
      sub301_1460 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1469_inst
    process(conv236_1301, conv238_1228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv236_1301, conv238_1228, tmp_var);
      sub310_1470 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1979_inst
    process(conv470_1866, conv454_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv470_1866, conv454_1742, tmp_var);
      sub518_1980 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1989_inst
    process(conv452_1815, conv454_1742) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv452_1815, conv454_1742, tmp_var);
      sub527_1990 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2513_inst
    process(conv692_2406, conv676_2283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv692_2406, conv676_2283, tmp_var);
      sub739_2514 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2523_inst
    process(conv674_2355, conv676_2283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv674_2355, conv676_2283, tmp_var);
      sub748_2524 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3039_inst
    process(conv909_2926, conv892_2796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv909_2926, conv892_2796, tmp_var);
      sub957_3040 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3049_inst
    process(conv890_2869, conv892_2796) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv890_2869, conv892_2796, tmp_var);
      sub966_3050 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3585_inst
    process(conv1133_3478, conv1116_3349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1133_3478, conv1116_3349, tmp_var);
      sub1180_3586 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3595_inst
    process(conv1114_3421, conv1116_3349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1114_3421, conv1116_3349, tmp_var);
      sub1189_3596 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4111_inst
    process(conv1350_3998, conv1335_3880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1350_3998, conv1335_3880, tmp_var);
      sub1398_4112 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4121_inst
    process(conv1333_3953, conv1335_3880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1333_3953, conv1335_3880, tmp_var);
      sub1407_4122 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4639_inst
    process(conv1571_4532, conv1556_4415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1571_4532, conv1556_4415, tmp_var);
      sub1618_4640 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4649_inst
    process(conv1554_4487, conv1556_4415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1554_4487, conv1556_4415, tmp_var);
      sub1627_4650 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_938_inst
    process(conv50_824, conv38_698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv50_824, conv38_698, tmp_var);
      sub_939 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_948_inst
    process(conv36_773, conv38_698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv36_773, conv38_698, tmp_var);
      sub99_949 <= tmp_var; --
    end process;
    -- shared split operator group (348) : array_obj_ref_1003_index_offset 
    ApIntAdd_group_348: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom120_1002_scaled;
      array_obj_ref_1003_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1003_index_offset_req_0;
      array_obj_ref_1003_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1003_index_offset_req_1;
      array_obj_ref_1003_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_348_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_348_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_348",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 348
    -- shared split operator group (349) : array_obj_ref_1028_index_offset 
    ApIntAdd_group_349: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom125_1027_scaled;
      array_obj_ref_1028_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1028_index_offset_req_0;
      array_obj_ref_1028_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1028_index_offset_req_1;
      array_obj_ref_1028_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_349_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_349_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_349",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 349
    -- shared split operator group (350) : array_obj_ref_1441_index_offset 
    ApIntAdd_group_350: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom288_1440_scaled;
      array_obj_ref_1441_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1441_index_offset_req_0;
      array_obj_ref_1441_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1441_index_offset_req_1;
      array_obj_ref_1441_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_350_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_350_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_350",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 350
    -- shared split operator group (351) : array_obj_ref_1524_index_offset 
    ApIntAdd_group_351: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom331_1523_scaled;
      array_obj_ref_1524_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1524_index_offset_req_0;
      array_obj_ref_1524_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1524_index_offset_req_1;
      array_obj_ref_1524_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_351_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_351_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_351",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 351
    -- shared split operator group (352) : array_obj_ref_1549_index_offset 
    ApIntAdd_group_352: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom336_1548_scaled;
      array_obj_ref_1549_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1549_index_offset_req_0;
      array_obj_ref_1549_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1549_index_offset_req_1;
      array_obj_ref_1549_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_352_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_352_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_352",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 352
    -- shared split operator group (353) : array_obj_ref_1961_index_offset 
    ApIntAdd_group_353: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom505_1960_scaled;
      array_obj_ref_1961_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1961_index_offset_req_0;
      array_obj_ref_1961_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1961_index_offset_req_1;
      array_obj_ref_1961_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_353_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_353_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_353",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 353
    -- shared split operator group (354) : array_obj_ref_2044_index_offset 
    ApIntAdd_group_354: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom548_2043_scaled;
      array_obj_ref_2044_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2044_index_offset_req_0;
      array_obj_ref_2044_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2044_index_offset_req_1;
      array_obj_ref_2044_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_354_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_354_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_354",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 354
    -- shared split operator group (355) : array_obj_ref_2069_index_offset 
    ApIntAdd_group_355: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom553_2068_scaled;
      array_obj_ref_2069_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2069_index_offset_req_0;
      array_obj_ref_2069_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2069_index_offset_req_1;
      array_obj_ref_2069_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_355_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_355_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_355",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 355
    -- shared split operator group (356) : array_obj_ref_2495_index_offset 
    ApIntAdd_group_356: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom726_2494_scaled;
      array_obj_ref_2495_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2495_index_offset_req_0;
      array_obj_ref_2495_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2495_index_offset_req_1;
      array_obj_ref_2495_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_356_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_356_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_356",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 356
    -- shared split operator group (357) : array_obj_ref_2578_index_offset 
    ApIntAdd_group_357: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom769_2577_scaled;
      array_obj_ref_2578_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2578_index_offset_req_0;
      array_obj_ref_2578_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2578_index_offset_req_1;
      array_obj_ref_2578_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_357_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_357_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_357",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 357
    -- shared split operator group (358) : array_obj_ref_2603_index_offset 
    ApIntAdd_group_358: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom774_2602_scaled;
      array_obj_ref_2603_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2603_index_offset_req_0;
      array_obj_ref_2603_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2603_index_offset_req_1;
      array_obj_ref_2603_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_358_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_358_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_358",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 358
    -- shared split operator group (359) : array_obj_ref_3021_index_offset 
    ApIntAdd_group_359: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom944_3020_scaled;
      array_obj_ref_3021_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3021_index_offset_req_0;
      array_obj_ref_3021_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3021_index_offset_req_1;
      array_obj_ref_3021_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_359_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_359_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_359",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 359
    -- shared split operator group (360) : array_obj_ref_3104_index_offset 
    ApIntAdd_group_360: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom987_3103_scaled;
      array_obj_ref_3104_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3104_index_offset_req_0;
      array_obj_ref_3104_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3104_index_offset_req_1;
      array_obj_ref_3104_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_360_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_360_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_360",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 360
    -- shared split operator group (361) : array_obj_ref_3129_index_offset 
    ApIntAdd_group_361: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom992_3128_scaled;
      array_obj_ref_3129_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3129_index_offset_req_0;
      array_obj_ref_3129_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3129_index_offset_req_1;
      array_obj_ref_3129_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_361_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_361_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_361",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 361
    -- shared split operator group (362) : array_obj_ref_3567_index_offset 
    ApIntAdd_group_362: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1167_3566_scaled;
      array_obj_ref_3567_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3567_index_offset_req_0;
      array_obj_ref_3567_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3567_index_offset_req_1;
      array_obj_ref_3567_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_362_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_362_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_362",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 362
    -- shared split operator group (363) : array_obj_ref_3650_index_offset 
    ApIntAdd_group_363: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1210_3649_scaled;
      array_obj_ref_3650_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3650_index_offset_req_0;
      array_obj_ref_3650_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3650_index_offset_req_1;
      array_obj_ref_3650_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_363_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_363_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_363",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 363
    -- shared split operator group (364) : array_obj_ref_3675_index_offset 
    ApIntAdd_group_364: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1215_3674_scaled;
      array_obj_ref_3675_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3675_index_offset_req_0;
      array_obj_ref_3675_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3675_index_offset_req_1;
      array_obj_ref_3675_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_364_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_364_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_364",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 364
    -- shared split operator group (365) : array_obj_ref_4093_index_offset 
    ApIntAdd_group_365: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1385_4092_scaled;
      array_obj_ref_4093_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4093_index_offset_req_0;
      array_obj_ref_4093_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4093_index_offset_req_1;
      array_obj_ref_4093_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_365_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_365_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_365",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 365
    -- shared split operator group (366) : array_obj_ref_4176_index_offset 
    ApIntAdd_group_366: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1428_4175_scaled;
      array_obj_ref_4176_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4176_index_offset_req_0;
      array_obj_ref_4176_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4176_index_offset_req_1;
      array_obj_ref_4176_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_366_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_366_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_366",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 366
    -- shared split operator group (367) : array_obj_ref_4201_index_offset 
    ApIntAdd_group_367: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1433_4200_scaled;
      array_obj_ref_4201_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4201_index_offset_req_0;
      array_obj_ref_4201_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4201_index_offset_req_1;
      array_obj_ref_4201_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_367_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_367_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_367",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 367
    -- shared split operator group (368) : array_obj_ref_4621_index_offset 
    ApIntAdd_group_368: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1605_4620_scaled;
      array_obj_ref_4621_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4621_index_offset_req_0;
      array_obj_ref_4621_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4621_index_offset_req_1;
      array_obj_ref_4621_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_368_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_368_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_368",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 368
    -- shared split operator group (369) : array_obj_ref_4704_index_offset 
    ApIntAdd_group_369: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1648_4703_scaled;
      array_obj_ref_4704_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4704_index_offset_req_0;
      array_obj_ref_4704_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4704_index_offset_req_1;
      array_obj_ref_4704_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_369_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_369_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_369",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 369
    -- shared split operator group (370) : array_obj_ref_4729_index_offset 
    ApIntAdd_group_370: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1653_4728_scaled;
      array_obj_ref_4729_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4729_index_offset_req_0;
      array_obj_ref_4729_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4729_index_offset_req_1;
      array_obj_ref_4729_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_370_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_370_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_370",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 370
    -- shared split operator group (371) : array_obj_ref_920_index_offset 
    ApIntAdd_group_371: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_919_scaled;
      array_obj_ref_920_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_920_index_offset_req_0;
      array_obj_ref_920_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_920_index_offset_req_1;
      array_obj_ref_920_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_371_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_371_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_371",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 371
    -- unary operator type_cast_1021_inst
    process(shr124_1018) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr124_1018, tmp_var);
      type_cast_1021_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1039_inst
    process(kx_x1_761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_761, tmp_var);
      type_cast_1039_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1078_inst
    process(inc_1075) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1075, tmp_var);
      type_cast_1078_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1122_inst
    process(inc155x_xix_x2_1112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc155x_xix_x2_1112, tmp_var);
      type_cast_1122_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1299_inst
    process(i184x_x2_1282) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i184x_x2_1282, tmp_var);
      type_cast_1299_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1350_inst
    process(j230x_x1_1276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j230x_x1_1276, tmp_var);
      type_cast_1350_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1395_inst
    process(k176x_x1_1289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k176x_x1_1289, tmp_var);
      type_cast_1395_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1400_inst
    process(j230x_x1_1276) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j230x_x1_1276, tmp_var);
      type_cast_1400_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1434_inst
    process(shr287_1431) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr287_1431, tmp_var);
      type_cast_1434_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1453_inst
    process(k176x_x1_1289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k176x_x1_1289, tmp_var);
      type_cast_1453_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1517_inst
    process(shr330_1514) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr330_1514, tmp_var);
      type_cast_1517_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1542_inst
    process(shr335_1539) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr335_1539, tmp_var);
      type_cast_1542_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1560_inst
    process(k176x_x1_1289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k176x_x1_1289, tmp_var);
      type_cast_1560_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1599_inst
    process(inc355_1596) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc355_1596, tmp_var);
      type_cast_1599_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1636_inst
    process(inc369x_xi184x_x2_1627) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc369x_xi184x_x2_1627, tmp_var);
      type_cast_1636_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1813_inst
    process(i396x_x2_1797) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i396x_x2_1797, tmp_var);
      type_cast_1813_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1864_inst
    process(j446x_x1_1803) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j446x_x1_1803, tmp_var);
      type_cast_1864_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1915_inst
    process(k392x_x1_1790) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k392x_x1_1790, tmp_var);
      type_cast_1915_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1920_inst
    process(j446x_x1_1803) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j446x_x1_1803, tmp_var);
      type_cast_1920_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1954_inst
    process(shr504_1951) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr504_1951, tmp_var);
      type_cast_1954_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1973_inst
    process(k392x_x1_1790) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k392x_x1_1790, tmp_var);
      type_cast_1973_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2037_inst
    process(shr547_2034) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr547_2034, tmp_var);
      type_cast_2037_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2062_inst
    process(shr552_2059) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr552_2059, tmp_var);
      type_cast_2062_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2080_inst
    process(k392x_x1_1790) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k392x_x1_1790, tmp_var);
      type_cast_2080_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2119_inst
    process(inc572_2116) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc572_2116, tmp_var);
      type_cast_2119_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2163_inst
    process(inc587x_xi396x_x2_2153) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc587x_xi396x_x2_2153, tmp_var);
      type_cast_2163_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2353_inst
    process(i618x_x2_2338) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i618x_x2_2338, tmp_var);
      type_cast_2353_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2404_inst
    process(j668x_x1_2344) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j668x_x1_2344, tmp_var);
      type_cast_2404_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2449_inst
    process(k610x_x1_2331) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k610x_x1_2331, tmp_var);
      type_cast_2449_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2454_inst
    process(j668x_x1_2344) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j668x_x1_2344, tmp_var);
      type_cast_2454_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2488_inst
    process(shr725_2485) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr725_2485, tmp_var);
      type_cast_2488_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2507_inst
    process(k610x_x1_2331) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k610x_x1_2331, tmp_var);
      type_cast_2507_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2571_inst
    process(shr768_2568) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr768_2568, tmp_var);
      type_cast_2571_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2596_inst
    process(shr773_2593) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr773_2593, tmp_var);
      type_cast_2596_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2614_inst
    process(k610x_x1_2331) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k610x_x1_2331, tmp_var);
      type_cast_2614_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2653_inst
    process(inc793_2650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc793_2650, tmp_var);
      type_cast_2653_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2690_inst
    process(inc807x_xi618x_x2_2681) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc807x_xi618x_x2_2681, tmp_var);
      type_cast_2690_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2867_inst
    process(i834x_x2_2851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i834x_x2_2851, tmp_var);
      type_cast_2867_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2924_inst
    process(j884x_x1_2857) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j884x_x1_2857, tmp_var);
      type_cast_2924_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2975_inst
    process(k830x_x1_2844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k830x_x1_2844, tmp_var);
      type_cast_2975_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2980_inst
    process(j884x_x1_2857) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j884x_x1_2857, tmp_var);
      type_cast_2980_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3014_inst
    process(shr943_3011) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr943_3011, tmp_var);
      type_cast_3014_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3033_inst
    process(k830x_x1_2844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k830x_x1_2844, tmp_var);
      type_cast_3033_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3097_inst
    process(shr986_3094) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr986_3094, tmp_var);
      type_cast_3097_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3122_inst
    process(shr991_3119) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr991_3119, tmp_var);
      type_cast_3122_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3140_inst
    process(k830x_x1_2844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k830x_x1_2844, tmp_var);
      type_cast_3140_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3179_inst
    process(inc1011_3176) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1011_3176, tmp_var);
      type_cast_3179_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3223_inst
    process(inc1026x_xi834x_x2_3213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1026x_xi834x_x2_3213, tmp_var);
      type_cast_3223_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3419_inst
    process(i1058x_x2_3404) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1058x_x2_3404, tmp_var);
      type_cast_3419_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3476_inst
    process(j1108x_x1_3410) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1108x_x1_3410, tmp_var);
      type_cast_3476_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3521_inst
    process(k1050x_x1_3397) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1050x_x1_3397, tmp_var);
      type_cast_3521_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3526_inst
    process(j1108x_x1_3410) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1108x_x1_3410, tmp_var);
      type_cast_3526_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3560_inst
    process(shr1166_3557) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1166_3557, tmp_var);
      type_cast_3560_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3579_inst
    process(k1050x_x1_3397) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1050x_x1_3397, tmp_var);
      type_cast_3579_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3643_inst
    process(shr1209_3640) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1209_3640, tmp_var);
      type_cast_3643_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3668_inst
    process(shr1214_3665) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1214_3665, tmp_var);
      type_cast_3668_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3686_inst
    process(k1050x_x1_3397) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1050x_x1_3397, tmp_var);
      type_cast_3686_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3725_inst
    process(inc1234_3722) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1234_3722, tmp_var);
      type_cast_3725_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3762_inst
    process(inc1248x_xi1058x_x2_3753) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1248x_xi1058x_x2_3753, tmp_var);
      type_cast_3762_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3951_inst
    process(i1276x_x2_3935) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1276x_x2_3935, tmp_var);
      type_cast_3951_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3996_inst
    process(j1327x_x1_3941) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1327x_x1_3941, tmp_var);
      type_cast_3996_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4047_inst
    process(k1272x_x1_3928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1272x_x1_3928, tmp_var);
      type_cast_4047_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4052_inst
    process(j1327x_x1_3941) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1327x_x1_3941, tmp_var);
      type_cast_4052_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4086_inst
    process(shr1384_4083) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1384_4083, tmp_var);
      type_cast_4086_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4105_inst
    process(k1272x_x1_3928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1272x_x1_3928, tmp_var);
      type_cast_4105_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4169_inst
    process(shr1427_4166) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1427_4166, tmp_var);
      type_cast_4169_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4194_inst
    process(shr1432_4191) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1432_4191, tmp_var);
      type_cast_4194_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4212_inst
    process(k1272x_x1_3928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1272x_x1_3928, tmp_var);
      type_cast_4212_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4251_inst
    process(inc1452_4248) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1452_4248, tmp_var);
      type_cast_4251_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4295_inst
    process(inc1467x_xi1276x_x2_4285) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1467x_xi1276x_x2_4285, tmp_var);
      type_cast_4295_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4485_inst
    process(i1497x_x2_4470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1497x_x2_4470, tmp_var);
      type_cast_4485_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4530_inst
    process(j1548x_x1_4476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1548x_x1_4476, tmp_var);
      type_cast_4530_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4575_inst
    process(k1489x_x1_4463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1489x_x1_4463, tmp_var);
      type_cast_4575_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4580_inst
    process(j1548x_x1_4476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1548x_x1_4476, tmp_var);
      type_cast_4580_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4614_inst
    process(shr1604_4611) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1604_4611, tmp_var);
      type_cast_4614_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4633_inst
    process(k1489x_x1_4463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1489x_x1_4463, tmp_var);
      type_cast_4633_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4697_inst
    process(shr1647_4694) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1647_4694, tmp_var);
      type_cast_4697_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4722_inst
    process(shr1652_4719) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1652_4719, tmp_var);
      type_cast_4722_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4740_inst
    process(k1489x_x1_4463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1489x_x1_4463, tmp_var);
      type_cast_4740_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4779_inst
    process(inc1672_4776) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1672_4776, tmp_var);
      type_cast_4779_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4816_inst
    process(inc1686x_xi1497x_x2_4807) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1686x_xi1497x_x2_4807, tmp_var);
      type_cast_4816_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_771_inst
    process(ix_x2_754) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_754, tmp_var);
      type_cast_771_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_822_inst
    process(jx_x1_747) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_747, tmp_var);
      type_cast_822_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_873_inst
    process(kx_x1_761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_761, tmp_var);
      type_cast_873_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_878_inst
    process(jx_x1_747) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_747, tmp_var);
      type_cast_878_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_913_inst
    process(shr_909) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_909, tmp_var);
      type_cast_913_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_932_inst
    process(kx_x1_761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_761, tmp_var);
      type_cast_932_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_996_inst
    process(shr119_993) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr119_993, tmp_var);
      type_cast_996_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_col_high_2657_load_0 LOAD_col_high_1882_load_0 LOAD_col_high_666_load_0 LOAD_col_high_840_load_0 LOAD_col_high_1082_load_0 LOAD_col_high_2942_load_0 LOAD_col_high_1368_load_0 LOAD_col_high_1603_load_0 LOAD_col_high_2123_load_0 LOAD_col_high_3729_load_0 LOAD_col_high_4014_load_0 LOAD_col_high_2422_load_0 LOAD_col_high_3183_load_0 LOAD_col_high_3494_load_0 LOAD_col_high_4255_load_0 LOAD_col_high_4783_load_0 LOAD_col_high_4548_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(16 downto 0);
      signal data_out: std_logic_vector(135 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 16 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 16 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 16 downto 0);
      signal guard_vector : std_logic_vector( 16 downto 0);
      constant inBUFs : IntegerArray(16 downto 0) := (16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(16 downto 0) := (16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(16 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false);
      constant guardBuffering: IntegerArray(16 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2);
      -- 
    begin -- 
      reqL_unguarded(16) <= LOAD_col_high_2657_load_0_req_0;
      reqL_unguarded(15) <= LOAD_col_high_1882_load_0_req_0;
      reqL_unguarded(14) <= LOAD_col_high_666_load_0_req_0;
      reqL_unguarded(13) <= LOAD_col_high_840_load_0_req_0;
      reqL_unguarded(12) <= LOAD_col_high_1082_load_0_req_0;
      reqL_unguarded(11) <= LOAD_col_high_2942_load_0_req_0;
      reqL_unguarded(10) <= LOAD_col_high_1368_load_0_req_0;
      reqL_unguarded(9) <= LOAD_col_high_1603_load_0_req_0;
      reqL_unguarded(8) <= LOAD_col_high_2123_load_0_req_0;
      reqL_unguarded(7) <= LOAD_col_high_3729_load_0_req_0;
      reqL_unguarded(6) <= LOAD_col_high_4014_load_0_req_0;
      reqL_unguarded(5) <= LOAD_col_high_2422_load_0_req_0;
      reqL_unguarded(4) <= LOAD_col_high_3183_load_0_req_0;
      reqL_unguarded(3) <= LOAD_col_high_3494_load_0_req_0;
      reqL_unguarded(2) <= LOAD_col_high_4255_load_0_req_0;
      reqL_unguarded(1) <= LOAD_col_high_4783_load_0_req_0;
      reqL_unguarded(0) <= LOAD_col_high_4548_load_0_req_0;
      LOAD_col_high_2657_load_0_ack_0 <= ackL_unguarded(16);
      LOAD_col_high_1882_load_0_ack_0 <= ackL_unguarded(15);
      LOAD_col_high_666_load_0_ack_0 <= ackL_unguarded(14);
      LOAD_col_high_840_load_0_ack_0 <= ackL_unguarded(13);
      LOAD_col_high_1082_load_0_ack_0 <= ackL_unguarded(12);
      LOAD_col_high_2942_load_0_ack_0 <= ackL_unguarded(11);
      LOAD_col_high_1368_load_0_ack_0 <= ackL_unguarded(10);
      LOAD_col_high_1603_load_0_ack_0 <= ackL_unguarded(9);
      LOAD_col_high_2123_load_0_ack_0 <= ackL_unguarded(8);
      LOAD_col_high_3729_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_col_high_4014_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_col_high_2422_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_col_high_3183_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_col_high_3494_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_col_high_4255_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_col_high_4783_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_col_high_4548_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(16) <= LOAD_col_high_2657_load_0_req_1;
      reqR_unguarded(15) <= LOAD_col_high_1882_load_0_req_1;
      reqR_unguarded(14) <= LOAD_col_high_666_load_0_req_1;
      reqR_unguarded(13) <= LOAD_col_high_840_load_0_req_1;
      reqR_unguarded(12) <= LOAD_col_high_1082_load_0_req_1;
      reqR_unguarded(11) <= LOAD_col_high_2942_load_0_req_1;
      reqR_unguarded(10) <= LOAD_col_high_1368_load_0_req_1;
      reqR_unguarded(9) <= LOAD_col_high_1603_load_0_req_1;
      reqR_unguarded(8) <= LOAD_col_high_2123_load_0_req_1;
      reqR_unguarded(7) <= LOAD_col_high_3729_load_0_req_1;
      reqR_unguarded(6) <= LOAD_col_high_4014_load_0_req_1;
      reqR_unguarded(5) <= LOAD_col_high_2422_load_0_req_1;
      reqR_unguarded(4) <= LOAD_col_high_3183_load_0_req_1;
      reqR_unguarded(3) <= LOAD_col_high_3494_load_0_req_1;
      reqR_unguarded(2) <= LOAD_col_high_4255_load_0_req_1;
      reqR_unguarded(1) <= LOAD_col_high_4783_load_0_req_1;
      reqR_unguarded(0) <= LOAD_col_high_4548_load_0_req_1;
      LOAD_col_high_2657_load_0_ack_1 <= ackR_unguarded(16);
      LOAD_col_high_1882_load_0_ack_1 <= ackR_unguarded(15);
      LOAD_col_high_666_load_0_ack_1 <= ackR_unguarded(14);
      LOAD_col_high_840_load_0_ack_1 <= ackR_unguarded(13);
      LOAD_col_high_1082_load_0_ack_1 <= ackR_unguarded(12);
      LOAD_col_high_2942_load_0_ack_1 <= ackR_unguarded(11);
      LOAD_col_high_1368_load_0_ack_1 <= ackR_unguarded(10);
      LOAD_col_high_1603_load_0_ack_1 <= ackR_unguarded(9);
      LOAD_col_high_2123_load_0_ack_1 <= ackR_unguarded(8);
      LOAD_col_high_3729_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_col_high_4014_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_col_high_2422_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_col_high_3183_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_col_high_3494_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_col_high_4255_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_col_high_4783_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_col_high_4548_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_16: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_16", num_slots => 1) -- 
        port map (req => reqL_unregulated(16), -- 
          ack => ackL_unregulated(16),
          regulated_req => reqL(16),
          regulated_ack => ackL(16),
          release_req => reqR(16),
          release_ack => ackR(16),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 17, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_col_high_2657_word_address_0 & LOAD_col_high_1882_word_address_0 & LOAD_col_high_666_word_address_0 & LOAD_col_high_840_word_address_0 & LOAD_col_high_1082_word_address_0 & LOAD_col_high_2942_word_address_0 & LOAD_col_high_1368_word_address_0 & LOAD_col_high_1603_word_address_0 & LOAD_col_high_2123_word_address_0 & LOAD_col_high_3729_word_address_0 & LOAD_col_high_4014_word_address_0 & LOAD_col_high_2422_word_address_0 & LOAD_col_high_3183_word_address_0 & LOAD_col_high_3494_word_address_0 & LOAD_col_high_4255_word_address_0 & LOAD_col_high_4783_word_address_0 & LOAD_col_high_4548_word_address_0;
      LOAD_col_high_2657_data_0 <= data_out(135 downto 128);
      LOAD_col_high_1882_data_0 <= data_out(127 downto 120);
      LOAD_col_high_666_data_0 <= data_out(119 downto 112);
      LOAD_col_high_840_data_0 <= data_out(111 downto 104);
      LOAD_col_high_1082_data_0 <= data_out(103 downto 96);
      LOAD_col_high_2942_data_0 <= data_out(95 downto 88);
      LOAD_col_high_1368_data_0 <= data_out(87 downto 80);
      LOAD_col_high_1603_data_0 <= data_out(79 downto 72);
      LOAD_col_high_2123_data_0 <= data_out(71 downto 64);
      LOAD_col_high_3729_data_0 <= data_out(63 downto 56);
      LOAD_col_high_4014_data_0 <= data_out(55 downto 48);
      LOAD_col_high_2422_data_0 <= data_out(47 downto 40);
      LOAD_col_high_3183_data_0 <= data_out(39 downto 32);
      LOAD_col_high_3494_data_0 <= data_out(31 downto 24);
      LOAD_col_high_4255_data_0 <= data_out(23 downto 16);
      LOAD_col_high_4783_data_0 <= data_out(15 downto 8);
      LOAD_col_high_4548_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 17,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 17,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : LOAD_depth_high_1714_load_0 LOAD_depth_high_663_load_0 LOAD_depth_high_1200_load_0 LOAD_depth_high_2768_load_0 LOAD_depth_high_2255_load_0 LOAD_depth_high_3852_load_0 LOAD_depth_high_3321_load_0 LOAD_depth_high_4387_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_depth_high_1714_load_0_req_0;
      reqL_unguarded(6) <= LOAD_depth_high_663_load_0_req_0;
      reqL_unguarded(5) <= LOAD_depth_high_1200_load_0_req_0;
      reqL_unguarded(4) <= LOAD_depth_high_2768_load_0_req_0;
      reqL_unguarded(3) <= LOAD_depth_high_2255_load_0_req_0;
      reqL_unguarded(2) <= LOAD_depth_high_3852_load_0_req_0;
      reqL_unguarded(1) <= LOAD_depth_high_3321_load_0_req_0;
      reqL_unguarded(0) <= LOAD_depth_high_4387_load_0_req_0;
      LOAD_depth_high_1714_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_depth_high_663_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_depth_high_1200_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_depth_high_2768_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_depth_high_2255_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_depth_high_3852_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_depth_high_3321_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_depth_high_4387_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_depth_high_1714_load_0_req_1;
      reqR_unguarded(6) <= LOAD_depth_high_663_load_0_req_1;
      reqR_unguarded(5) <= LOAD_depth_high_1200_load_0_req_1;
      reqR_unguarded(4) <= LOAD_depth_high_2768_load_0_req_1;
      reqR_unguarded(3) <= LOAD_depth_high_2255_load_0_req_1;
      reqR_unguarded(2) <= LOAD_depth_high_3852_load_0_req_1;
      reqR_unguarded(1) <= LOAD_depth_high_3321_load_0_req_1;
      reqR_unguarded(0) <= LOAD_depth_high_4387_load_0_req_1;
      LOAD_depth_high_1714_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_depth_high_663_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_depth_high_1200_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_depth_high_2768_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_depth_high_2255_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_depth_high_3852_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_depth_high_3321_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_depth_high_4387_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_depth_high_1714_word_address_0 & LOAD_depth_high_663_word_address_0 & LOAD_depth_high_1200_word_address_0 & LOAD_depth_high_2768_word_address_0 & LOAD_depth_high_2255_word_address_0 & LOAD_depth_high_3852_word_address_0 & LOAD_depth_high_3321_word_address_0 & LOAD_depth_high_4387_word_address_0;
      LOAD_depth_high_1714_data_0 <= data_out(63 downto 56);
      LOAD_depth_high_663_data_0 <= data_out(55 downto 48);
      LOAD_depth_high_1200_data_0 <= data_out(47 downto 40);
      LOAD_depth_high_2768_data_0 <= data_out(39 downto 32);
      LOAD_depth_high_2255_data_0 <= data_out(31 downto 24);
      LOAD_depth_high_3852_data_0 <= data_out(23 downto 16);
      LOAD_depth_high_3321_data_0 <= data_out(15 downto 8);
      LOAD_depth_high_4387_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(7 downto 0),
          mtag => memory_space_4_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : LOAD_out_col_high_1720_load_0 LOAD_out_col_high_672_load_0 LOAD_out_col_high_3858_load_0 LOAD_out_col_high_1206_load_0 LOAD_out_col_high_2774_load_0 LOAD_out_col_high_2261_load_0 LOAD_out_col_high_3327_load_0 LOAD_out_col_high_4393_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_out_col_high_1720_load_0_req_0;
      reqL_unguarded(6) <= LOAD_out_col_high_672_load_0_req_0;
      reqL_unguarded(5) <= LOAD_out_col_high_3858_load_0_req_0;
      reqL_unguarded(4) <= LOAD_out_col_high_1206_load_0_req_0;
      reqL_unguarded(3) <= LOAD_out_col_high_2774_load_0_req_0;
      reqL_unguarded(2) <= LOAD_out_col_high_2261_load_0_req_0;
      reqL_unguarded(1) <= LOAD_out_col_high_3327_load_0_req_0;
      reqL_unguarded(0) <= LOAD_out_col_high_4393_load_0_req_0;
      LOAD_out_col_high_1720_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_out_col_high_672_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_out_col_high_3858_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_out_col_high_1206_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_out_col_high_2774_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_out_col_high_2261_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_out_col_high_3327_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_out_col_high_4393_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_out_col_high_1720_load_0_req_1;
      reqR_unguarded(6) <= LOAD_out_col_high_672_load_0_req_1;
      reqR_unguarded(5) <= LOAD_out_col_high_3858_load_0_req_1;
      reqR_unguarded(4) <= LOAD_out_col_high_1206_load_0_req_1;
      reqR_unguarded(3) <= LOAD_out_col_high_2774_load_0_req_1;
      reqR_unguarded(2) <= LOAD_out_col_high_2261_load_0_req_1;
      reqR_unguarded(1) <= LOAD_out_col_high_3327_load_0_req_1;
      reqR_unguarded(0) <= LOAD_out_col_high_4393_load_0_req_1;
      LOAD_out_col_high_1720_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_out_col_high_672_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_out_col_high_3858_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_out_col_high_1206_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_out_col_high_2774_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_out_col_high_2261_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_out_col_high_3327_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_out_col_high_4393_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_out_col_high_1720_word_address_0 & LOAD_out_col_high_672_word_address_0 & LOAD_out_col_high_3858_word_address_0 & LOAD_out_col_high_1206_word_address_0 & LOAD_out_col_high_2774_word_address_0 & LOAD_out_col_high_2261_word_address_0 & LOAD_out_col_high_3327_word_address_0 & LOAD_out_col_high_4393_word_address_0;
      LOAD_out_col_high_1720_data_0 <= data_out(63 downto 56);
      LOAD_out_col_high_672_data_0 <= data_out(55 downto 48);
      LOAD_out_col_high_3858_data_0 <= data_out(47 downto 40);
      LOAD_out_col_high_1206_data_0 <= data_out(39 downto 32);
      LOAD_out_col_high_2774_data_0 <= data_out(31 downto 24);
      LOAD_out_col_high_2261_data_0 <= data_out(23 downto 16);
      LOAD_out_col_high_3327_data_0 <= data_out(15 downto 8);
      LOAD_out_col_high_4393_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(7 downto 0),
          mtag => memory_space_6_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : LOAD_out_depth_high_1717_load_0 LOAD_out_depth_high_669_load_0 LOAD_out_depth_high_1203_load_0 LOAD_out_depth_high_2771_load_0 LOAD_out_depth_high_3855_load_0 LOAD_out_depth_high_2258_load_0 LOAD_out_depth_high_3324_load_0 LOAD_out_depth_high_4390_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_out_depth_high_1717_load_0_req_0;
      reqL_unguarded(6) <= LOAD_out_depth_high_669_load_0_req_0;
      reqL_unguarded(5) <= LOAD_out_depth_high_1203_load_0_req_0;
      reqL_unguarded(4) <= LOAD_out_depth_high_2771_load_0_req_0;
      reqL_unguarded(3) <= LOAD_out_depth_high_3855_load_0_req_0;
      reqL_unguarded(2) <= LOAD_out_depth_high_2258_load_0_req_0;
      reqL_unguarded(1) <= LOAD_out_depth_high_3324_load_0_req_0;
      reqL_unguarded(0) <= LOAD_out_depth_high_4390_load_0_req_0;
      LOAD_out_depth_high_1717_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_out_depth_high_669_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_out_depth_high_1203_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_out_depth_high_2771_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_out_depth_high_3855_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_out_depth_high_2258_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_out_depth_high_3324_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_out_depth_high_4390_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_out_depth_high_1717_load_0_req_1;
      reqR_unguarded(6) <= LOAD_out_depth_high_669_load_0_req_1;
      reqR_unguarded(5) <= LOAD_out_depth_high_1203_load_0_req_1;
      reqR_unguarded(4) <= LOAD_out_depth_high_2771_load_0_req_1;
      reqR_unguarded(3) <= LOAD_out_depth_high_3855_load_0_req_1;
      reqR_unguarded(2) <= LOAD_out_depth_high_2258_load_0_req_1;
      reqR_unguarded(1) <= LOAD_out_depth_high_3324_load_0_req_1;
      reqR_unguarded(0) <= LOAD_out_depth_high_4390_load_0_req_1;
      LOAD_out_depth_high_1717_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_out_depth_high_669_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_out_depth_high_1203_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_out_depth_high_2771_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_out_depth_high_3855_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_out_depth_high_2258_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_out_depth_high_3324_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_out_depth_high_4390_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_out_depth_high_1717_word_address_0 & LOAD_out_depth_high_669_word_address_0 & LOAD_out_depth_high_1203_word_address_0 & LOAD_out_depth_high_2771_word_address_0 & LOAD_out_depth_high_3855_word_address_0 & LOAD_out_depth_high_2258_word_address_0 & LOAD_out_depth_high_3324_word_address_0 & LOAD_out_depth_high_4390_word_address_0;
      LOAD_out_depth_high_1717_data_0 <= data_out(63 downto 56);
      LOAD_out_depth_high_669_data_0 <= data_out(55 downto 48);
      LOAD_out_depth_high_1203_data_0 <= data_out(47 downto 40);
      LOAD_out_depth_high_2771_data_0 <= data_out(39 downto 32);
      LOAD_out_depth_high_3855_data_0 <= data_out(31 downto 24);
      LOAD_out_depth_high_2258_data_0 <= data_out(23 downto 16);
      LOAD_out_depth_high_3324_data_0 <= data_out(15 downto 8);
      LOAD_out_depth_high_4390_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : LOAD_pad_1711_load_0 LOAD_pad_660_load_0 LOAD_pad_1197_load_0 LOAD_pad_2765_load_0 LOAD_pad_2252_load_0 LOAD_pad_3849_load_0 LOAD_pad_3318_load_0 LOAD_pad_4384_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_pad_1711_load_0_req_0;
      reqL_unguarded(6) <= LOAD_pad_660_load_0_req_0;
      reqL_unguarded(5) <= LOAD_pad_1197_load_0_req_0;
      reqL_unguarded(4) <= LOAD_pad_2765_load_0_req_0;
      reqL_unguarded(3) <= LOAD_pad_2252_load_0_req_0;
      reqL_unguarded(2) <= LOAD_pad_3849_load_0_req_0;
      reqL_unguarded(1) <= LOAD_pad_3318_load_0_req_0;
      reqL_unguarded(0) <= LOAD_pad_4384_load_0_req_0;
      LOAD_pad_1711_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_pad_660_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_pad_1197_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_pad_2765_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_pad_2252_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_pad_3849_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_pad_3318_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_pad_4384_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_pad_1711_load_0_req_1;
      reqR_unguarded(6) <= LOAD_pad_660_load_0_req_1;
      reqR_unguarded(5) <= LOAD_pad_1197_load_0_req_1;
      reqR_unguarded(4) <= LOAD_pad_2765_load_0_req_1;
      reqR_unguarded(3) <= LOAD_pad_2252_load_0_req_1;
      reqR_unguarded(2) <= LOAD_pad_3849_load_0_req_1;
      reqR_unguarded(1) <= LOAD_pad_3318_load_0_req_1;
      reqR_unguarded(0) <= LOAD_pad_4384_load_0_req_1;
      LOAD_pad_1711_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_pad_660_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_pad_1197_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_pad_2765_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_pad_2252_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_pad_3849_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_pad_3318_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_pad_4384_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_1711_word_address_0 & LOAD_pad_660_word_address_0 & LOAD_pad_1197_word_address_0 & LOAD_pad_2765_word_address_0 & LOAD_pad_2252_word_address_0 & LOAD_pad_3849_word_address_0 & LOAD_pad_3318_word_address_0 & LOAD_pad_4384_word_address_0;
      LOAD_pad_1711_data_0 <= data_out(63 downto 56);
      LOAD_pad_660_data_0 <= data_out(55 downto 48);
      LOAD_pad_1197_data_0 <= data_out(47 downto 40);
      LOAD_pad_2765_data_0 <= data_out(39 downto 32);
      LOAD_pad_2252_data_0 <= data_out(31 downto 24);
      LOAD_pad_3849_data_0 <= data_out(23 downto 16);
      LOAD_pad_3318_data_0 <= data_out(15 downto 8);
      LOAD_pad_4384_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_9_lr_req(0),
          mack => memory_space_9_lr_ack(0),
          maddr => memory_space_9_lr_addr(0 downto 0),
          mtag => memory_space_9_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_9_lc_req(0),
          mack => memory_space_9_lc_ack(0),
          mdata => memory_space_9_lc_data(7 downto 0),
          mtag => memory_space_9_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : LOAD_row_high_789_load_0 LOAD_row_high_1831_load_0 LOAD_row_high_2885_load_0 LOAD_row_high_1126_load_0 LOAD_row_high_2694_load_0 LOAD_row_high_1317_load_0 LOAD_row_high_1640_load_0 LOAD_row_high_2167_load_0 LOAD_row_high_3766_load_0 LOAD_row_high_3969_load_0 LOAD_row_high_2371_load_0 LOAD_row_high_4820_load_0 LOAD_row_high_3227_load_0 LOAD_row_high_3437_load_0 LOAD_row_high_4299_load_0 LOAD_row_high_4503_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= LOAD_row_high_789_load_0_req_0;
      reqL_unguarded(14) <= LOAD_row_high_1831_load_0_req_0;
      reqL_unguarded(13) <= LOAD_row_high_2885_load_0_req_0;
      reqL_unguarded(12) <= LOAD_row_high_1126_load_0_req_0;
      reqL_unguarded(11) <= LOAD_row_high_2694_load_0_req_0;
      reqL_unguarded(10) <= LOAD_row_high_1317_load_0_req_0;
      reqL_unguarded(9) <= LOAD_row_high_1640_load_0_req_0;
      reqL_unguarded(8) <= LOAD_row_high_2167_load_0_req_0;
      reqL_unguarded(7) <= LOAD_row_high_3766_load_0_req_0;
      reqL_unguarded(6) <= LOAD_row_high_3969_load_0_req_0;
      reqL_unguarded(5) <= LOAD_row_high_2371_load_0_req_0;
      reqL_unguarded(4) <= LOAD_row_high_4820_load_0_req_0;
      reqL_unguarded(3) <= LOAD_row_high_3227_load_0_req_0;
      reqL_unguarded(2) <= LOAD_row_high_3437_load_0_req_0;
      reqL_unguarded(1) <= LOAD_row_high_4299_load_0_req_0;
      reqL_unguarded(0) <= LOAD_row_high_4503_load_0_req_0;
      LOAD_row_high_789_load_0_ack_0 <= ackL_unguarded(15);
      LOAD_row_high_1831_load_0_ack_0 <= ackL_unguarded(14);
      LOAD_row_high_2885_load_0_ack_0 <= ackL_unguarded(13);
      LOAD_row_high_1126_load_0_ack_0 <= ackL_unguarded(12);
      LOAD_row_high_2694_load_0_ack_0 <= ackL_unguarded(11);
      LOAD_row_high_1317_load_0_ack_0 <= ackL_unguarded(10);
      LOAD_row_high_1640_load_0_ack_0 <= ackL_unguarded(9);
      LOAD_row_high_2167_load_0_ack_0 <= ackL_unguarded(8);
      LOAD_row_high_3766_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_row_high_3969_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_row_high_2371_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_row_high_4820_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_row_high_3227_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_row_high_3437_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_row_high_4299_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_row_high_4503_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= LOAD_row_high_789_load_0_req_1;
      reqR_unguarded(14) <= LOAD_row_high_1831_load_0_req_1;
      reqR_unguarded(13) <= LOAD_row_high_2885_load_0_req_1;
      reqR_unguarded(12) <= LOAD_row_high_1126_load_0_req_1;
      reqR_unguarded(11) <= LOAD_row_high_2694_load_0_req_1;
      reqR_unguarded(10) <= LOAD_row_high_1317_load_0_req_1;
      reqR_unguarded(9) <= LOAD_row_high_1640_load_0_req_1;
      reqR_unguarded(8) <= LOAD_row_high_2167_load_0_req_1;
      reqR_unguarded(7) <= LOAD_row_high_3766_load_0_req_1;
      reqR_unguarded(6) <= LOAD_row_high_3969_load_0_req_1;
      reqR_unguarded(5) <= LOAD_row_high_2371_load_0_req_1;
      reqR_unguarded(4) <= LOAD_row_high_4820_load_0_req_1;
      reqR_unguarded(3) <= LOAD_row_high_3227_load_0_req_1;
      reqR_unguarded(2) <= LOAD_row_high_3437_load_0_req_1;
      reqR_unguarded(1) <= LOAD_row_high_4299_load_0_req_1;
      reqR_unguarded(0) <= LOAD_row_high_4503_load_0_req_1;
      LOAD_row_high_789_load_0_ack_1 <= ackR_unguarded(15);
      LOAD_row_high_1831_load_0_ack_1 <= ackR_unguarded(14);
      LOAD_row_high_2885_load_0_ack_1 <= ackR_unguarded(13);
      LOAD_row_high_1126_load_0_ack_1 <= ackR_unguarded(12);
      LOAD_row_high_2694_load_0_ack_1 <= ackR_unguarded(11);
      LOAD_row_high_1317_load_0_ack_1 <= ackR_unguarded(10);
      LOAD_row_high_1640_load_0_ack_1 <= ackR_unguarded(9);
      LOAD_row_high_2167_load_0_ack_1 <= ackR_unguarded(8);
      LOAD_row_high_3766_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_row_high_3969_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_row_high_2371_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_row_high_4820_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_row_high_3227_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_row_high_3437_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_row_high_4299_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_row_high_4503_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      LoadGroup5_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_row_high_789_word_address_0 & LOAD_row_high_1831_word_address_0 & LOAD_row_high_2885_word_address_0 & LOAD_row_high_1126_word_address_0 & LOAD_row_high_2694_word_address_0 & LOAD_row_high_1317_word_address_0 & LOAD_row_high_1640_word_address_0 & LOAD_row_high_2167_word_address_0 & LOAD_row_high_3766_word_address_0 & LOAD_row_high_3969_word_address_0 & LOAD_row_high_2371_word_address_0 & LOAD_row_high_4820_word_address_0 & LOAD_row_high_3227_word_address_0 & LOAD_row_high_3437_word_address_0 & LOAD_row_high_4299_word_address_0 & LOAD_row_high_4503_word_address_0;
      LOAD_row_high_789_data_0 <= data_out(127 downto 120);
      LOAD_row_high_1831_data_0 <= data_out(119 downto 112);
      LOAD_row_high_2885_data_0 <= data_out(111 downto 104);
      LOAD_row_high_1126_data_0 <= data_out(103 downto 96);
      LOAD_row_high_2694_data_0 <= data_out(95 downto 88);
      LOAD_row_high_1317_data_0 <= data_out(87 downto 80);
      LOAD_row_high_1640_data_0 <= data_out(79 downto 72);
      LOAD_row_high_2167_data_0 <= data_out(71 downto 64);
      LOAD_row_high_3766_data_0 <= data_out(63 downto 56);
      LOAD_row_high_3969_data_0 <= data_out(55 downto 48);
      LOAD_row_high_2371_data_0 <= data_out(47 downto 40);
      LOAD_row_high_4820_data_0 <= data_out(39 downto 32);
      LOAD_row_high_3227_data_0 <= data_out(31 downto 24);
      LOAD_row_high_3437_data_0 <= data_out(23 downto 16);
      LOAD_row_high_4299_data_0 <= data_out(15 downto 8);
      LOAD_row_high_4503_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 1,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(0),
          mack => memory_space_10_lr_ack(0),
          maddr => memory_space_10_lr_addr(0 downto 0),
          mtag => memory_space_10_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 8,
        num_reqs => 16,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(0),
          mack => memory_space_10_lc_ack(0),
          mdata => memory_space_10_lc_data(7 downto 0),
          mtag => memory_space_10_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_1008_load_0 ptr_deref_2583_load_0 ptr_deref_1529_load_0 ptr_deref_2049_load_0 ptr_deref_3655_load_0 ptr_deref_3109_load_0 ptr_deref_4181_load_0 ptr_deref_4709_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= ptr_deref_1008_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_2583_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_1529_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_2049_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_3655_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_3109_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_4181_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4709_load_0_req_0;
      ptr_deref_1008_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_2583_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_1529_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_2049_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_3655_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_3109_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_4181_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4709_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_1008_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_2583_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_1529_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_2049_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_3655_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_3109_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_4181_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4709_load_0_req_1;
      ptr_deref_1008_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_2583_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_1529_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_2049_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_3655_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_3109_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_4181_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4709_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup6_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1008_word_address_0 & ptr_deref_2583_word_address_0 & ptr_deref_1529_word_address_0 & ptr_deref_2049_word_address_0 & ptr_deref_3655_word_address_0 & ptr_deref_3109_word_address_0 & ptr_deref_4181_word_address_0 & ptr_deref_4709_word_address_0;
      ptr_deref_1008_data_0 <= data_out(511 downto 448);
      ptr_deref_2583_data_0 <= data_out(447 downto 384);
      ptr_deref_1529_data_0 <= data_out(383 downto 320);
      ptr_deref_2049_data_0 <= data_out(319 downto 256);
      ptr_deref_3655_data_0 <= data_out(255 downto 192);
      ptr_deref_3109_data_0 <= data_out(191 downto 128);
      ptr_deref_4181_data_0 <= data_out(127 downto 64);
      ptr_deref_4709_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 14,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 64,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared store operator group (0) : ptr_deref_2607_store_0 ptr_deref_1965_store_0 ptr_deref_2499_store_0 ptr_deref_924_store_0 ptr_deref_1032_store_0 ptr_deref_1445_store_0 ptr_deref_1553_store_0 ptr_deref_3025_store_0 ptr_deref_3571_store_0 ptr_deref_2073_store_0 ptr_deref_4097_store_0 ptr_deref_3133_store_0 ptr_deref_4625_store_0 ptr_deref_3679_store_0 ptr_deref_4733_store_0 ptr_deref_4205_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(223 downto 0);
      signal data_in: std_logic_vector(1023 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_2607_store_0_req_0;
      reqL_unguarded(14) <= ptr_deref_1965_store_0_req_0;
      reqL_unguarded(13) <= ptr_deref_2499_store_0_req_0;
      reqL_unguarded(12) <= ptr_deref_924_store_0_req_0;
      reqL_unguarded(11) <= ptr_deref_1032_store_0_req_0;
      reqL_unguarded(10) <= ptr_deref_1445_store_0_req_0;
      reqL_unguarded(9) <= ptr_deref_1553_store_0_req_0;
      reqL_unguarded(8) <= ptr_deref_3025_store_0_req_0;
      reqL_unguarded(7) <= ptr_deref_3571_store_0_req_0;
      reqL_unguarded(6) <= ptr_deref_2073_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_4097_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_3133_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_4625_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_3679_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_4733_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4205_store_0_req_0;
      ptr_deref_2607_store_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_1965_store_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_2499_store_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_924_store_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_1032_store_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_1445_store_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_1553_store_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_3025_store_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_3571_store_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_2073_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_4097_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_3133_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_4625_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_3679_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_4733_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4205_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_2607_store_0_req_1;
      reqR_unguarded(14) <= ptr_deref_1965_store_0_req_1;
      reqR_unguarded(13) <= ptr_deref_2499_store_0_req_1;
      reqR_unguarded(12) <= ptr_deref_924_store_0_req_1;
      reqR_unguarded(11) <= ptr_deref_1032_store_0_req_1;
      reqR_unguarded(10) <= ptr_deref_1445_store_0_req_1;
      reqR_unguarded(9) <= ptr_deref_1553_store_0_req_1;
      reqR_unguarded(8) <= ptr_deref_3025_store_0_req_1;
      reqR_unguarded(7) <= ptr_deref_3571_store_0_req_1;
      reqR_unguarded(6) <= ptr_deref_2073_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_4097_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_3133_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_4625_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_3679_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_4733_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4205_store_0_req_1;
      ptr_deref_2607_store_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_1965_store_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_2499_store_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_924_store_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_1032_store_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_1445_store_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_1553_store_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_3025_store_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_3571_store_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_2073_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_4097_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_3133_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_4625_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_3679_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_4733_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4205_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_11: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_12: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_13: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_14: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_15: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2607_word_address_0 & ptr_deref_1965_word_address_0 & ptr_deref_2499_word_address_0 & ptr_deref_924_word_address_0 & ptr_deref_1032_word_address_0 & ptr_deref_1445_word_address_0 & ptr_deref_1553_word_address_0 & ptr_deref_3025_word_address_0 & ptr_deref_3571_word_address_0 & ptr_deref_2073_word_address_0 & ptr_deref_4097_word_address_0 & ptr_deref_3133_word_address_0 & ptr_deref_4625_word_address_0 & ptr_deref_3679_word_address_0 & ptr_deref_4733_word_address_0 & ptr_deref_4205_word_address_0;
      data_in <= ptr_deref_2607_data_0 & ptr_deref_1965_data_0 & ptr_deref_2499_data_0 & ptr_deref_924_data_0 & ptr_deref_1032_data_0 & ptr_deref_1445_data_0 & ptr_deref_1553_data_0 & ptr_deref_3025_data_0 & ptr_deref_3571_data_0 & ptr_deref_2073_data_0 & ptr_deref_4097_data_0 & ptr_deref_3133_data_0 & ptr_deref_4625_data_0 & ptr_deref_3679_data_0 & ptr_deref_4733_data_0 & ptr_deref_4205_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 16,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared call operator group (0) : call_stmt_4866_call 
    sendOutput_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_4866_call_req_0;
      call_stmt_4866_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_4866_call_req_1;
      call_stmt_4866_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_0_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_657_call 
    testConfigure_call_group_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_657_call_req_0;
      call_stmt_657_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_657_call_req_1;
      call_stmt_657_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_1_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_657 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_10
  signal memory_space_10_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_10_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_10_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_10_lr_tag : std_logic_vector(43 downto 0);
  signal memory_space_10_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_10_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_10_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_10_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_10_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_10_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_10_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(43 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_3
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(41 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(41 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(41 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_9
  signal memory_space_9_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_9_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_9_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_9_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_9_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_9_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_10_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_9_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_9_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_10_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_9_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_9_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_9_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_9_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_9_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_9_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_10_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_10_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_10_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_10_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(21 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(4 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(1 downto 1),
      memory_space_6_lr_tag => memory_space_6_lr_tag(41 downto 21),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(15 downto 8),
      memory_space_6_lc_tag => memory_space_6_lc_tag(7 downto 4),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(41 downto 21),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 8),
      memory_space_7_lc_tag => memory_space_7_lc_tag(7 downto 4),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(0 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(17 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(7 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(0 downto 0),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(1 downto 1),
      memory_space_2_lr_tag => memory_space_2_lr_tag(43 downto 22),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(15 downto 8),
      memory_space_2_lc_tag => memory_space_2_lc_tag(9 downto 5),
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(1 downto 1),
      memory_space_4_lr_tag => memory_space_4_lr_tag(41 downto 21),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(15 downto 8),
      memory_space_4_lc_tag => memory_space_4_lc_tag(7 downto 4),
      memory_space_10_lr_req => memory_space_10_lr_req(1 downto 1),
      memory_space_10_lr_ack => memory_space_10_lr_ack(1 downto 1),
      memory_space_10_lr_addr => memory_space_10_lr_addr(1 downto 1),
      memory_space_10_lr_tag => memory_space_10_lr_tag(43 downto 22),
      memory_space_10_lc_req => memory_space_10_lc_req(1 downto 1),
      memory_space_10_lc_ack => memory_space_10_lc_ack(1 downto 1),
      memory_space_10_lc_data => memory_space_10_lc_data(15 downto 8),
      memory_space_10_lc_tag => memory_space_10_lc_tag(9 downto 5),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(7 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(21 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(0 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(7 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(20 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(3 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(6 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(31 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(1 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(1 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(0 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(7 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(20 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(3 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(7 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(20 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(3 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(7 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(17 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(0 downto 0),
      memory_space_9_sr_req => memory_space_9_sr_req(0 downto 0),
      memory_space_9_sr_ack => memory_space_9_sr_ack(0 downto 0),
      memory_space_9_sr_addr => memory_space_9_sr_addr(0 downto 0),
      memory_space_9_sr_data => memory_space_9_sr_data(7 downto 0),
      memory_space_9_sr_tag => memory_space_9_sr_tag(20 downto 0),
      memory_space_9_sc_req => memory_space_9_sc_req(0 downto 0),
      memory_space_9_sc_ack => memory_space_9_sc_ack(0 downto 0),
      memory_space_9_sc_tag => memory_space_9_sc_tag(3 downto 0),
      memory_space_10_sr_req => memory_space_10_sr_req(0 downto 0),
      memory_space_10_sr_ack => memory_space_10_sr_ack(0 downto 0),
      memory_space_10_sr_addr => memory_space_10_sr_addr(0 downto 0),
      memory_space_10_sr_data => memory_space_10_sr_data(7 downto 0),
      memory_space_10_sr_tag => memory_space_10_sr_tag(21 downto 0),
      memory_space_10_sc_req => memory_space_10_sc_req(0 downto 0),
      memory_space_10_sc_ack => memory_space_10_sc_ack(0 downto 0),
      memory_space_10_sc_tag => memory_space_10_sc_tag(4 downto 0),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(21 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(7 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(4 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(0 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(20 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(7 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(0 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(20 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(7 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(3 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(20 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(7 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 0),
      memory_space_9_lr_req => memory_space_9_lr_req(0 downto 0),
      memory_space_9_lr_ack => memory_space_9_lr_ack(0 downto 0),
      memory_space_9_lr_addr => memory_space_9_lr_addr(0 downto 0),
      memory_space_9_lr_tag => memory_space_9_lr_tag(20 downto 0),
      memory_space_9_lc_req => memory_space_9_lc_req(0 downto 0),
      memory_space_9_lc_ack => memory_space_9_lc_ack(0 downto 0),
      memory_space_9_lc_data => memory_space_9_lc_data(7 downto 0),
      memory_space_9_lc_tag => memory_space_9_lc_tag(3 downto 0),
      memory_space_10_lr_req => memory_space_10_lr_req(0 downto 0),
      memory_space_10_lr_ack => memory_space_10_lr_ack(0 downto 0),
      memory_space_10_lr_addr => memory_space_10_lr_addr(0 downto 0),
      memory_space_10_lr_tag => memory_space_10_lr_tag(21 downto 0),
      memory_space_10_lc_req => memory_space_10_lc_req(0 downto 0),
      memory_space_10_lc_ack => memory_space_10_lc_ack(0 downto 0),
      memory_space_10_lc_data => memory_space_10_lc_data(7 downto 0),
      memory_space_10_lc_tag => memory_space_10_lc_tag(4 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(21 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(4 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_10: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_10",
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_10_lr_addr,
      lr_req_in => memory_space_10_lr_req,
      lr_ack_out => memory_space_10_lr_ack,
      lr_tag_in => memory_space_10_lr_tag,
      lc_req_in => memory_space_10_lc_req,
      lc_ack_out => memory_space_10_lc_ack,
      lc_data_out => memory_space_10_lc_data,
      lc_tag_out => memory_space_10_lc_tag,
      sr_addr_in => memory_space_10_sr_addr,
      sr_data_in => memory_space_10_sr_data,
      sr_req_in => memory_space_10_sr_req,
      sr_ack_out => memory_space_10_sr_ack,
      sr_tag_in => memory_space_10_sr_tag,
      sc_req_in=> memory_space_10_sc_req,
      sc_ack_out => memory_space_10_sc_ack,
      sc_tag_out => memory_space_10_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_5: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_9: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_9",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_9_lr_addr,
      lr_req_in => memory_space_9_lr_req,
      lr_ack_out => memory_space_9_lr_ack,
      lr_tag_in => memory_space_9_lr_tag,
      lc_req_in => memory_space_9_lc_req,
      lc_ack_out => memory_space_9_lc_ack,
      lc_data_out => memory_space_9_lc_data,
      lc_tag_out => memory_space_9_lc_tag,
      sr_addr_in => memory_space_9_sr_addr,
      sr_data_in => memory_space_9_sr_data,
      sr_req_in => memory_space_9_sr_req,
      sr_ack_out => memory_space_9_sr_ack,
      sr_tag_in => memory_space_9_sr_tag,
      sc_req_in=> memory_space_9_sc_req,
      sc_ack_out => memory_space_9_sc_ack,
      sc_tag_out => memory_space_9_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
